#
# Copyright (C) 2003 Taiwan Semiconductor Manufacturing Company, Ltd.
# Confidential Information of TSMC, Ltd.
# Use subject to TSMC Design Service Division license.
# 
# Library : tcbn90g 
# File    : tcbn90g_9lm.lef
# Date    : Mon Dec 29 18:46:28 2003
#-------------------------------------------------------------------------
# 
# Routing layer capacitance definition issues
# ===========================================
#
#     In LEF file, two keywords are used by Silicon Ensemble to calculate
#
#   routing capacitance, i.e., CAPACITANCE CPRESQDIST and EDGECAPACITANCE,
#
#   where CAPACITANCE CPRESQDIST and EDGECAPACITANCE are used to calculate
#
#   area and fringe capacitance of each routing segment, respectively.
#
#
#
#      For deep sub-micron process, coupling capacitance plays a major role
#
#   in determining a net's total capacitance. For TSMC 0.35um 1P4M process,
#
#   a minimum width metal 4 wire with two other metal 4 wires run in
#
#   parallel with minimum spacing, its coupling capacitance is greater 80%
#
#   of the total capacitance. This percentage will drop to ~ 30% if the
#
#   other two parallel metal 4 wires are 5 times minimum spacing away.
#
#   (Please refer to TSMC 0.35um 1P4M SPICE Documents.) It is clear that
#
#   routing wire's capacitance greatly depends on its neighboring wires.
#
#   Unfortunately, there is no parameter in LEF to describe this effect.
#
#
#
#      To compensate coupling effect in LEF, as suggested in Cadence "
#
#   Timing-Driven Design Flow Guide" (Product version 5.1, page 3-11, May
#
#   29,1998), coupling values should be added to EDGECAPACITANCE. However,
#
#   only one value can be used. If the coupling capacitance with minimum
#
#   spacing is used, the extracted capacitance will be too larger for
#
#   non-minimum spacing wires. If another value is selected, it will also
#
#   make other patterns capacitance in-accurate.
#
#
#
#      For TSMC released LEF files, several test cases are used to calibrate
#
#   EDGECAPACITANCE values in LEF, where EDGECAPACITANCE is defined as the
#
#   sum of fringe capacitance and coupling capacitance of a metal wire with
#
#   two parallel wires at 2*minimum spacing away. For our test cases, the
#
#   mean difference of the extracted capacitance by using LEF file and using
#
#   Coeffgen (SE built-in field solver) is about 15%.~20% . Please note
#
#   that, as mentioned earlier, the capacitance compensation for LEF is
#
#   allowed for only one patterns. Usually, the majority one is used and it
#
#   is case dependent. Therefore, our result may be different case by case.
#
#   However, user can easily adjust the value of EDGECAPACITANCE for his
#
#   specific design by using the method described in Cadence "Timing-Driven
#
#   Design Flow Guide" or using our method described above.
#
#
#
#      In Silicon Ensemble, capacitance data defined in LEF files are used
#
#   to speed up routing process. More accurate RC extractors should be used
#
#   for final verification.
#
#-------------------------------------------------------------------------

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  CAPACITANCE PICOFARADS 10 ;
  CURRENT MILLIAMPS 10000 ;
  VOLTAGE VOLTS 1000 ;
  FREQUENCY MEGAHERTZ 10 ;
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;


LAYER PO
  TYPE MASTERSLICE ;
END PO


LAYER CO
  TYPE CUT ;
END CO


LAYER M1
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET 0 ;
  WIDTH .12 ;
  DIRECTION HORIZONTAL ;
  EDGECAPACITANCE 6.17E-05 ;
  RESISTANCE RPERSQ 1.05E-01 ;
  CAPACITANCE CPERSQDIST 1.091667E-04 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;


  WIREEXTENSION 0.11 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.12    0.12    0.12    0.12
  WIDTH    0.18         0.12    0.17    0.17    0.17
  WIDTH    1.50         0.12    0.17    0.50    0.50
  WIDTH    4.50         0.12    0.17    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.18 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  AREA 0.058 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.250000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.12 1.0 12 ;
    TABLEENTRIES
              3.536  34.648  423.557 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.12 1 ;
    TABLEENTRIES 
              0.2 1.96 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.12 0.24 0.5 1 5 12 ;
    TABLEENTRIES  
              2.325 3.786 6.544 11.523 50.183 117.556 ;
END M1


LAYER VIA1
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA1


LAYER M2
  TYPE ROUTING ;
  PITCH .32 ;
  OFFSET .16 ;
  WIDTH .14 ;
  DIRECTION VERTICAL ;
  THICKNESS .325 ;
  EDGECAPACITANCE 5.83E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M2


LAYER VIA2
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA2


LAYER M3
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET 0 ;
  WIDTH .14 ;
  DIRECTION HORIZONTAL ;
  THICKNESS .325 ;
  EDGECAPACITANCE 5.83E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;


  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50 
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M3


LAYER VIA3
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA3


LAYER M4
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET .16 ;
  WIDTH .14 ;
  DIRECTION VERTICAL ;
  THICKNESS .325 ;
  EDGECAPACITANCE 5.83E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M4


LAYER VIA4
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA4


LAYER M5
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET 0 ;
  WIDTH .14 ;
  DIRECTION HORIZONTAL ;

  THICKNESS .325 ;

  EDGECAPACITANCE 5.83E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50 
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ; 
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M5


LAYER VIA5
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA5


LAYER M6
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET .16 ;
  WIDTH .14 ;
  DIRECTION VERTICAL ;
  THICKNESS .325 ;
  EDGECAPACITANCE 5.83E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M6


LAYER VIA6
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.17 ADJACENTCUTS 3 WITHIN 0.19 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.093 ;
END VIA6


LAYER M7
  TYPE ROUTING ;
  PITCH .28 ;
  OFFSET 0 ;
  WIDTH .14 ;
  DIRECTION HORIZONTAL ;

  THICKNESS .325 ;
  EDGECAPACITANCE 5.93E-05 ;
  RESISTANCE RPERSQ 7.8E-02 ;
  CAPACITANCE CPERSQDIST 9.71429E-05 ;

  MINIMUMCUT 2 WIDTH 0.42 ;
  MINIMUMCUT 4 WIDTH 0.98 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.98 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.70 LENGTH 0.70 WITHIN 1.0 ;
  MINIMUMCUT 2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.0 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.115 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    0.52    1.50    4.50
  WIDTH    0.00         0.14    0.14    0.14    0.14
  WIDTH    0.21         0.14    0.19    0.19    0.19
  WIDTH    1.50         0.14    0.19    0.50    0.50
  WIDTH    4.50         0.14    0.19    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50 
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.07 ;
  MINENCLOSEDAREA 0.20 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.21 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.325000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.14 1.0 12 ;
    TABLEENTRIES
              2.758  22.521 275.312 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.14 1 ;
    TABLEENTRIES 
              0.312 2.548 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.14 0.28 0.56 1 5 12 ;
    TABLEENTRIES  
              1.660 2.656 4.375 6.894 28.857 67.024 ;

END M7


LAYER VIA7
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.713 ;
END VIA7


LAYER M8
  TYPE ROUTING ;
  PITCH .84 ;
  OFFSET .16 ;
  WIDTH .42 ;
  DIRECTION VERTICAL ;
  EDGECAPACITANCE 1.3309E-04 ;
  RESISTANCE RPERSQ 2.5E-02 ;
  CAPACITANCE CPERSQDIST 5.78571E-05 ;

  MINIMUMCUT 2 WIDTH 1.80 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.26 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    1.50    4.50
  WIDTH    0.00         0.42    0.42    0.42
  WIDTH    1.50         0.42    0.50    0.50
  WIDTH    4.50         0.42    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.565 ;
  MINENCLOSEDAREA 0.565 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.42 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.900000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 43027 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.42 1.0 12 ;
    TABLEENTRIES
              17.819  43.657 533.682 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.42 1 ;
    TABLEENTRIES 
              2.880 7.056 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.42 0.63 0.84 1 5 12 ;
    TABLEENTRIES  
              4.833 6.090 7.201 7.986 23.532 47.948 ;

END M8


LAYER VIA8
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;

  AntennaAreaRatio 20.000000 ;
  AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.059 20 ) ( 0.060 912 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;

  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    TABLEENTRIES 
              0.713 ;
END VIA8


LAYER M9
  TYPE ROUTING ;
  PITCH .84 ;
  OFFSET 0 ;
  WIDTH .42 ;
  DIRECTION HORIZONTAL ;
  EDGECAPACITANCE 7.58E-05 ;
  RESISTANCE RPERSQ 2.5E-02 ;
  CAPACITANCE CPERSQDIST 5.78571E-05 ;

  EDGECAPACITANCE .67E-04 ;
  RESISTANCE RPERSQ .25E-01 ;
  CAPACITANCE CPERSQDIST .58E-04 ;

  MINIMUMCUT 2 WIDTH 1.80 ;
  MINIMUMCUT 2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;

  WIREEXTENSION 0.26 ;
  MAXWIDTH 12.0 ;
  SPACINGTABLE
  PARALLELRUNLENGTH     0.00    1.50    4.50
  WIDTH    0.00         0.42    0.42    0.42
  WIDTH    1.50         0.42    0.50    0.50
  WIDTH    4.50         0.42    0.50    1.50 ;

  SPACINGTABLE
  INFLUENCE
  WIDTH 1.50 WITHIN 0.50 SPACING 0.50
  WIDTH 4.50 WITHIN 1.50 SPACING 1.50 ;

  AREA 0.565 ;
  MINENCLOSEDAREA 0.565 ;
  MINENCLOSEDAREA 0.80 WIDTH 0.42 ;
  MINENCLOSEDAREA 3.20 WIDTH 1.50 ;
  MINENCLOSEDAREA 7.20 WIDTH 3.00 ;
  MINENCLOSEDAREA 20.2 WIDTH 4.50 ;
  MINENCLOSEDAREA 51.8 WIDTH 7.50 ;

  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 100 100 ;
  DENSITYCHECKSTEP 50 ;
  FILLACTIVESPACING 2.0 ;

  Thickness 0.900000 ;
  AntennaAreaRatio 500.000000 ;
  AntennaCumAreaRatio 5000.000000 ;
  AntennaCumDiffAreaRatio PWL ( ( 0 5000 ) ( 0.059 5000 ) ( 0.060 50480 ) ( 0.5 54000 ) ( 1 58000 ) ( 1.5 62000 ) ) ;

  ACCURRENTDENSITY PEAK 
    FREQUENCY 500 ;
    WIDTH     0.42 1.0 12 ;
    TABLEENTRIES
              17.819  43.657 533.682 ; 
  ACCURRENTDENSITY AVERAGE
    FREQUENCY 500 ;
    WIDTH     0.42 1 ;
    TABLEENTRIES 
              2.880 7.056 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 500 ;
    WIDTH     0.42 0.63 0.84 1 5 12 ;
    TABLEENTRIES  
              4.833 6.090 7.201 7.986 23.532 47.948 ;

END M9


LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP


VIA VIA12 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.115 -0.070 0.115 0.070 ;
  LAYER VIA1 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M2 ;
    RECT -0.115 -0.070 0.115 0.070 ;
END VIA12


VIA VIA12R90 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M1 ;
    RECT -0.070 -0.115 0.070 0.115 ;
  LAYER VIA1 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M2 ;
    RECT -0.070 -0.115 0.070 0.115 ;
END VIA12R90


VIA VIA12_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M1 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA1 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M2 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA12_DBLCUT_H


VIA VIA12_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M1 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA1 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M2 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA12_DBLCUT_V


VIA VIA12_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M1 ;
    RECT -0.255 -0.210  0.255  0.210 ;
  LAYER VIA1 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M2 ;
    RECT -0.210 -0.255  0.210  0.255 ; 
END VIA12_QUADCUT


VIA VIA23 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M2 ;
    RECT -0.070 -0.115 0.070 0.115 ;
  LAYER VIA2 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M3 ;
    RECT -0.115 -0.070 0.115 0.070 ;
END VIA23


VIA VIA23NORTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M2 ;
        RECT -0.070 -0.115 0.070 0.385 ;
    LAYER VIA2 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M3 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA23NORTH


VIA VIA23SOUTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M2 ;
        RECT -0.070 -0.385 0.070 0.115 ;
    LAYER VIA2 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M3 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA23SOUTH


VIA VIA23_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M2 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA2 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M3 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA23_DBLCUT_H


VIA VIA23_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M2 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA2 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M3 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA23_DBLCUT_V


VIA VIA23_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M2 ;     
    RECT -0.210 -0.255  0.210  0.255 ;
  LAYER VIA2 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M3 ;
    RECT -0.255 -0.210  0.255  0.210 ;
END VIA23_QUADCUT


VIA VIA34 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M3 ;
    RECT -0.115 -0.070 0.115 0.070 ;
  LAYER VIA3 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M4 ;
    RECT -0.070 -0.115 0.070 0.115 ;
END VIA34


VIA VIA34EAST DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M3 ;
        RECT -0.115 -0.070 0.385 0.070 ;
    LAYER VIA3 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M4 ;
        RECT -0.070 -0.115 0.070 0.115 ;
END VIA34EAST


VIA VIA34WEST DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M3 ;
        RECT -0.385 -0.070 0.115 0.070 ;
    LAYER VIA3 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M4 ;
        RECT -0.070 -0.115 0.070 0.115 ;
END VIA34WEST


VIA VIA34_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M3 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA3 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M4 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA34_DBLCUT_H


VIA VIA34_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M3 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA3 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M4 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA34_DBLCUT_V


VIA VIA34_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M3 ;
    RECT -0.255 -0.210  0.255  0.210 ;
  LAYER VIA3 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M4 ;
    RECT -0.210 -0.255  0.210  0.255 ;
END VIA34_QUADCUT


VIA VIA45 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M4 ;
    RECT -0.070 -0.115 0.070 0.115 ;
  LAYER VIA4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M5 ;
    RECT -0.115 -0.070 0.115 0.070 ;
END VIA45


VIA VIA45NORTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6000000000 ;
    LAYER M4 ;
        RECT -0.070 -0.115 0.070 0.385 ;
    LAYER VIA4 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M5 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA45NORTH


VIA VIA45SOUTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6000000000 ;
    LAYER M4 ;
        RECT -0.070 -0.385 0.070 0.115 ;
    LAYER VIA4 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M5 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA45SOUTH


VIA VIA45_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M4 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA4 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M5 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA45_DBLCUT_H


VIA VIA45_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M4 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA4 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M5 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA45_DBLCUT_V


VIA VIA45_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M4 ;
    RECT -0.210 -0.255  0.210  0.255 ;
  LAYER VIA4 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M5 ;
    RECT -0.255 -0.210  0.255  0.210 ;
END VIA45_QUADCUT


VIA VIA56 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M5 ;
    RECT -0.115 -0.070 0.115 0.070 ;
  LAYER VIA5 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M6 ;
    RECT -0.070 -0.115 0.070 0.115 ;
END VIA56


VIA VIA56EAST DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6000000000 ;
    LAYER M5 ;
        RECT -0.115 -0.070 0.385 0.070 ;
    LAYER VIA5 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M6 ;
        RECT -0.070 -0.115 0.070 0.115 ;
END VIA56EAST


VIA VIA56WEST DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6000000000 ;
    LAYER M5 ;
        RECT -0.385 -0.070 0.115 0.070 ;
    LAYER VIA5 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M6 ;
        RECT -0.070 -0.115 0.070 0.115 ;
END VIA56WEST


VIA VIA56_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M5 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA5 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M6 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA56_DBLCUT_H


VIA VIA56_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M5 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA5 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M6 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA56_DBLCUT_V


VIA VIA56_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M5 ;
    RECT -0.255 -0.210  0.255  0.210 ;
  LAYER VIA5 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M6 ;
    RECT -0.210 -0.255  0.210  0.255 ;
END VIA56_QUADCUT


VIA VIA67 DEFAULT
  RESISTANCE 1.6 ;
  LAYER M6 ;
    RECT -0.070 -0.115 0.070 0.115 ;
  LAYER VIA6 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M7 ;
    RECT -0.115 -0.070 0.115 0.070 ;
END VIA67


VIA VIA67NORTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M6 ;
        RECT -0.070 -0.115 0.070 0.385 ;
    LAYER VIA6 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M7 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA67NORTH


VIA VIA67SOUTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 1.6 ;
    LAYER M6 ;
        RECT -0.070 -0.385 0.070 0.115 ;
    LAYER VIA6 ;
        RECT -0.065 -0.065 0.065 0.065 ;
    LAYER M7 ;
        RECT -0.115 -0.070 0.115 0.070 ;
END VIA67SOUTH


VIA VIA67_DBLCUT_H DEFAULT
  RESISTANCE 0.8 ;
  LAYER M6 ;
    RECT -0.255 -0.070 0.255 0.070 ;
  LAYER VIA6 ;
    RECT -0.205 -0.065 -0.075 0.065 ;
    RECT  0.075 -0.065  0.205 0.065 ;
  LAYER M7 ;
    RECT -0.255 -0.070 0.255 0.070 ;
END VIA67_DBLCUT_H


VIA VIA67_DBLCUT_V DEFAULT
  RESISTANCE 0.8 ;
  LAYER M6 ;
    RECT -0.070 -0.255 0.070 0.255 ;
  LAYER VIA6 ;
    RECT -0.065 -0.205  0.065 -0.075 ;
    RECT -0.065  0.075  0.065 0.205 ;
  LAYER M7 ;
    RECT -0.070 -0.255 0.070 0.255 ;
END VIA67_DBLCUT_V


VIA VIA67_QUADCUT DEFAULT
  RESISTANCE 0.4 ;
  LAYER M6 ;
    RECT -0.210 -0.255  0.210  0.255 ;
  LAYER VIA6 ;
    RECT  0.075  0.075  0.205  0.205 ;
    RECT -0.205  0.075 -0.075  0.205 ;
    RECT -0.205 -0.205 -0.075 -0.075 ;
    RECT  0.075 -0.205  0.205 -0.075 ;
  LAYER M7 ;
    RECT -0.255 -0.210  0.255  0.210 ;
END VIA67_QUADCUT


VIA VIA78 DEFAULT
  RESISTANCE 0.45000000000 ;
  LAYER M7 ;
    RECT -0.260 -0.210 0.260 0.210 ;
  LAYER VIA7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M8 ;
    RECT -0.210 -0.210 0.210 0.210 ;
END VIA78


VIA VIA78R90 DEFAULT
  RESISTANCE 0.45 ;
  LAYER M7 ;
    RECT -0.210 -0.260 0.210 0.260 ;
  LAYER VIA7 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M8 ;
    RECT -0.210 -0.210 0.210 0.210 ;
END VIA78R90


VIA VIA78_DBLCUT_H DEFAULT
  RESISTANCE 0.225 ;
  LAYER M7 ;
    RECT -0.610 -0.210 0.610 0.210 ;
  LAYER VIA7 ;
    RECT -0.530 -0.180 -0.170 0.180 ;
    RECT  0.170 -0.180  0.530 0.180 ;
  LAYER M8 ;
    RECT -0.610 -0.210 0.610 0.210 ;
END VIA78_DBLCUT_H


VIA VIA78_DBLCUT_V DEFAULT
  RESISTANCE 0.225 ;
  LAYER M7 ;
    RECT -0.210 -0.610 0.210 0.610 ;
  LAYER VIA7 ;
    RECT -0.180 -0.530  0.180 -0.170 ;
    RECT -0.180  0.170  0.180  0.530 ;
  LAYER M8 ;
    RECT -0.210 -0.610 0.210 0.610 ;
END VIA78_DBLCUT_V


VIA VIA78_QUADCUT DEFAULT
  RESISTANCE 0.1125 ;
  LAYER M7 ;
    RECT -0.710 -0.660  0.710  0.660 ;
  LAYER VIA7 ;
    RECT  0.270  0.270  0.630  0.630 ;
    RECT -0.630  0.270 -0.270  0.630 ;
    RECT -0.630 -0.630 -0.270 -0.270 ;
    RECT  0.270 -0.630  0.630 -0.270 ;
  LAYER M8 ;
    RECT -0.660 -0.710  0.660  0.710 ;
END VIA78_QUADCUT


VIA VIA89 DEFAULT
  RESISTANCE 0.45000000000 ;
  LAYER M8 ;
    RECT -0.210 -0.210 0.210 0.210 ;
  LAYER VIA8 ;
    RECT -0.180 -0.180 0.180 0.180 ;
  LAYER M9 ;
    RECT -0.210 -0.210 0.210 0.210 ;
END VIA89


VIA VIA89NORTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.4500000000 ;
    LAYER M8 ;
        RECT -0.210 -0.260 0.210 1.090 ;
    LAYER VIA8 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER M9 ;
        RECT -0.260 -0.210 0.260 0.210 ;
END VIA89NORTH


VIA VIA89SOUTH DEFAULT TOPOFSTACKONLY
    RESISTANCE 0.4500000000 ;
    LAYER M8 ;
        RECT -0.210 -1.090 0.210 0.260 ;
    LAYER VIA8 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER M9 ;
        RECT -0.260 -0.210 0.260 0.210 ;
END VIA89SOUTH


VIA VIA89_DBLCUT_H DEFAULT
  RESISTANCE 0.225 ;
  LAYER M8 ;
    RECT -0.610 -0.210 0.610 0.210 ;
  LAYER VIA8 ;
    RECT -0.530 -0.180 -0.170 0.180 ;
    RECT  0.170 -0.180  0.530 0.180 ;
  LAYER M9 ;
    RECT -0.610 -0.210 0.610 0.210 ;
END VIA89_DBLCUT_H


VIA VIA89_DBLCUT_V DEFAULT
  RESISTANCE 0.225 ;
  LAYER M8 ;
    RECT -0.210 -0.610 0.210 0.610 ;
  LAYER VIA8 ;
    RECT -0.180 -0.530  0.180 -0.170 ;
    RECT -0.180  0.170  0.180  0.530 ;
  LAYER M9 ;
    RECT -0.210 -0.610 0.210 0.610 ;
END VIA89_DBLCUT_V


VIA VIA89_QUADCUT DEFAULT
  RESISTANCE 0.1125 ;
  LAYER M8 ;
    RECT -0.660 -0.710  0.660  0.710 ;
  LAYER VIA8 ;
    RECT  0.270  0.270  0.630  0.630 ;
    RECT -0.630  0.270 -0.270  0.630 ;
    RECT -0.630 -0.630 -0.270 -0.270 ;
    RECT  0.270 -0.630  0.630 -0.270 ;
  LAYER M9 ;
    RECT -0.710 -0.660  0.710  0.660 ;
END VIA89_QUADCUT


VIARULE VIAGEN12 GENERATE
   LAYER M1 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.12 TO 12.00 ;
   LAYER M2 ;
       ENCLOSURE .5E-01 .5E-02 ;
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA1 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ;
       SPACING .30 BY .30 ;    
END VIAGEN12        


VIARULE VIAGEN23 GENERATE
   LAYER M2 ;
       ENCLOSURE .5E-01 .5E-02 ;  
       WIDTH 0.14 TO 12.00 ;
   LAYER M3 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA2 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ; 
       SPACING .30 BY .30 ;    
END VIAGEN23


VIARULE VIAGEN34 GENERATE
   LAYER M3 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER M4 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA3 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ; 
       SPACING .30 BY .30 ;    
END VIAGEN34


VIARULE VIAGEN45 GENERATE
   LAYER M4 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER M5 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA4 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ; 
       SPACING .30 BY .30 ;    
END VIAGEN45


VIARULE VIAGEN56 GENERATE
   LAYER M5 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER M6 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA5 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ; 
       SPACING .30 BY .30 ;    
END VIAGEN56


VIARULE VIAGEN67 GENERATE
   LAYER M6 ;
       ENCLOSURE .5E-01 .5E-02  ;
       WIDTH 0.14 TO 12.00 ;
   LAYER M7 ;
       ENCLOSURE .5E-01 .5E-02 ; 
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA6 ;
       RECT -.65E-01 -.65E-01 .65E-01 .65E-01 ; 
       SPACING .30 BY .30 ;     
END VIAGEN67


VIARULE VIAGEN78 GENERATE
   LAYER M7 ;
       ENCLOSURE .8E-01 .3E-01  ;
       WIDTH 0.14 TO 12.00 ;
   LAYER M8 ;
       ENCLOSURE .8E-01 .3E-01  ;
       WIDTH 0.14 TO 12.00 ;
   LAYER VIA7 ;
       RECT -.18 -.18 .18 .18 ; 
       SPACING .90 BY .90 ;    
END VIAGEN78


VIARULE VIAGEN89 GENERATE
    LAYER M8 ;
       ENCLOSURE .8E-01 .3E-01  ;
       WIDTH 0.14 TO 12.00 ;
    LAYER M9 ;
       ENCLOSURE .8E-01 .3E-01  ;
       WIDTH 0.14 TO 12.00 ;
    LAYER VIA8 ;
       RECT -.18 -.18 .18 .18 ; 
       SPACING .90 BY .90 ;    
 END VIAGEN89           


MAXVIASTACK 4 RANGE M1 M7 ;


VIARULE TURN1 GENERATE
LAYER M1 ;
DIRECTION HORIZONTAL ;
LAYER M1 ;
DIRECTION VERTICAL ;
END TURN1


VIARULE TURN2 GENERATE
LAYER M2 ;
DIRECTION HORIZONTAL ;
LAYER M2 ;
DIRECTION VERTICAL ;
END TURN2


VIARULE TURN3 GENERATE
LAYER M3 ;
DIRECTION HORIZONTAL ;
LAYER M3 ;
DIRECTION VERTICAL ;
END TURN3


VIARULE TURN4 GENERATE
LAYER M4 ;
DIRECTION HORIZONTAL ;
LAYER M4 ;
DIRECTION VERTICAL ;
END TURN4


VIARULE TURN5 GENERATE
LAYER M5 ;
DIRECTION HORIZONTAL ;
LAYER M5 ;
DIRECTION VERTICAL ;
END TURN5


VIARULE TURN6 GENERATE
LAYER M6 ;
DIRECTION HORIZONTAL ;
LAYER M6 ;
DIRECTION VERTICAL ;
END TURN6


VIARULE TURN7 GENERATE
LAYER M7 ;
DIRECTION HORIZONTAL ;
LAYER M7 ;
DIRECTION VERTICAL ;
END TURN7


VIARULE TURN8 GENERATE
LAYER M8 ;
DIRECTION HORIZONTAL ;
LAYER M8 ;
DIRECTION VERTICAL ;
END TURN8


VIARULE TURN9 GENERATE
LAYER M9 ;
DIRECTION HORIZONTAL ;
LAYER M9 ;
DIRECTION VERTICAL ;
END TURN9


SPACING
  SAMENET VIA8 VIA8 .34 ;
  SAMENET VIA7 VIA7 .34 ;
  SAMENET VIA6 VIA6 .15 ;
  SAMENET VIA5 VIA5 .15 ;
  SAMENET VIA4 VIA4 .15 ;
  SAMENET VIA3 VIA3 .15 ;
  SAMENET VIA2 VIA2 .15 ;
  SAMENET VIA1 VIA1 .15 ;
  SAMENET VIA7 VIA8 0 STACK ;
  SAMENET VIA6 VIA7 0 STACK ;
  SAMENET VIA5 VIA6 0 STACK ;
  SAMENET VIA4 VIA5 0 STACK ;
  SAMENET VIA3 VIA4 0 STACK ;
  SAMENET VIA2 VIA3 0 STACK ;
  SAMENET VIA1 VIA2 0 STACK ;
  SAMENET M9 M9 .42 ;
  SAMENET M8 M8 .42 STACK ;
  SAMENET M7 M7 .14 STACK ;
  SAMENET M6 M6 .14 STACK ;
  SAMENET M5 M5 .14 STACK ;
  SAMENET M4 M4 .14 STACK ;
  SAMENET M3 M3 .14 STACK ;
  SAMENET M2 M2 .14 STACK ;
  SAMENET M1 M1 .12 ; 
END SPACING


SITE core
  SIZE .32 BY 2.52 ;
  CLASS CORE ;
  SYMMETRY Y  ;
END core



MACRO AN2D0
    CLASS CORE ;
    FOREIGN AN2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.910 1.040 2.100 ;
        RECT  1.030 0.420 1.040 0.610 ;
        RECT  1.040 0.420 1.190 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.265 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.600 0.300 ;
        RECT  0.600 -0.300 0.820 0.340 ;
        RECT  0.820 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.650 2.820 ;
        RECT  0.650 1.690 0.770 2.820 ;
        RECT  0.770 1.385 0.800 2.820 ;
        RECT  0.800 1.385 0.920 1.810 ;
        RECT  0.800 2.220 1.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.530 1.410 0.550 1.570 ;
        RECT  0.390 0.725 0.530 2.090 ;
        RECT  0.060 0.725 0.390 0.885 ;
        RECT  0.290 1.930 0.390 2.090 ;
    END
END AN2D0

MACRO AN2D1
    CLASS CORE ;
    FOREIGN AN2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.350 0.420 1.510 2.100 ;
        RECT  1.510 1.960 1.540 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.900 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.910 0.300 ;
        RECT  0.910 -0.300 1.130 0.340 ;
        RECT  1.130 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.910 2.820 ;
        RECT  0.910 2.180 1.130 2.820 ;
        RECT  1.130 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.710 1.230 1.800 ;
        RECT  0.220 0.710 1.070 0.870 ;
        RECT  0.470 1.640 1.070 1.800 ;
    END
END AN2D1

MACRO AN2D2
    CLASS CORE ;
    FOREIGN AN2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.960 1.310 2.100 ;
        RECT  1.310 1.390 1.370 2.100 ;
        RECT  1.310 0.420 1.370 0.900 ;
        RECT  1.370 0.420 1.470 2.100 ;
        RECT  1.470 1.960 1.500 2.100 ;
        RECT  1.470 0.780 1.510 1.515 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.870 0.300 ;
        RECT  0.870 -0.300 1.090 0.340 ;
        RECT  1.090 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.890 2.820 ;
        RECT  0.890 2.180 1.110 2.820 ;
        RECT  1.110 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.030 0.760 1.190 1.760 ;
        RECT  0.420 0.760 1.030 0.880 ;
        RECT  0.710 1.640 1.030 1.760 ;
        RECT  0.490 1.640 0.710 2.060 ;
        RECT  0.200 0.460 0.420 0.880 ;
    END
END AN2D2

MACRO AN2D4
    CLASS CORE ;
    FOREIGN AN2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.650 2.190 2.030 ;
        RECT  1.810 0.490 2.190 0.870 ;
        RECT  2.190 0.490 2.610 2.030 ;
        RECT  2.610 1.650 2.720 2.030 ;
        RECT  2.610 0.490 2.720 0.870 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.750 0.250 1.515 ;
        RECT  0.250 0.750 1.280 0.870 ;
        RECT  1.280 0.750 1.440 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.420 0.300 ;
        RECT  1.420 -0.300 1.640 0.340 ;
        RECT  1.640 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 1.080 1.900 1.240 ;
        RECT  1.570 0.470 1.690 1.510 ;
        RECT  0.750 0.470 1.570 0.630 ;
        RECT  1.310 1.390 1.570 1.510 ;
        RECT  1.310 1.960 1.340 2.100 ;
        RECT  1.150 1.390 1.310 2.100 ;
        RECT  0.610 1.390 1.150 1.510 ;
        RECT  1.120 1.960 1.150 2.100 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 1.390 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  1.810 0.490 1.975 0.870 ;
        RECT  1.810 1.650 1.975 2.030 ;
    END
END AN2D4

MACRO AN2D8
    CLASS CORE ;
    FOREIGN AN2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.640 3.470 2.020 ;
        RECT  2.500 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 4.950 2.020 ;
        RECT  3.890 0.500 4.950 0.880 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.030 1.235 ;
        RECT  1.030 0.760 1.190 1.235 ;
        RECT  1.190 0.760 1.970 0.880 ;
        RECT  1.970 0.760 2.130 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.030 0.490 1.510 ;
        RECT  0.490 1.390 1.370 1.510 ;
        RECT  1.370 1.005 1.490 1.510 ;
        RECT  1.490 1.005 1.830 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.820 0.300 ;
        RECT  0.820 -0.300 1.040 0.340 ;
        RECT  1.040 -0.300 2.100 0.300 ;
        RECT  2.100 -0.300 2.320 0.340 ;
        RECT  2.320 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.370 1.080 3.170 1.240 ;
        RECT  2.250 0.470 2.370 1.510 ;
        RECT  0.150 0.470 2.250 0.630 ;
        RECT  1.990 1.390 2.250 1.510 ;
        RECT  1.990 1.960 2.020 2.100 ;
        RECT  1.830 1.390 1.990 2.100 ;
        RECT  1.300 1.630 1.830 1.750 ;
        RECT  1.800 1.960 1.830 2.100 ;
        RECT  1.300 1.960 1.330 2.100 ;
        RECT  1.140 1.630 1.300 2.100 ;
        RECT  0.610 1.630 1.140 1.750 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 1.630 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  2.500 0.500 3.255 0.880 ;
        RECT  2.500 1.640 3.255 2.020 ;
        RECT  4.105 0.500 4.950 0.880 ;
        RECT  4.105 1.640 4.950 2.020 ;
    END
END AN2D8

MACRO AN3D0
    CLASS CORE ;
    FOREIGN AN3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.580 1.830 1.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.050 1.220 1.270 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.230 0.300 ;
        RECT  1.230 -0.300 1.450 0.340 ;
        RECT  1.450 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.630 1.550 1.820 ;
        RECT  0.290 0.630 1.390 0.790 ;
        RECT  0.070 1.660 1.390 1.820 ;
    END
END AN3D0

MACRO AN3D1
    CLASS CORE ;
    FOREIGN AN3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.670 0.420 1.830 2.100 ;
        RECT  1.830 1.960 1.860 2.100 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.970 1.210 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.130 0.300 ;
        RECT  1.130 -0.300 1.350 0.340 ;
        RECT  1.350 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.380 0.630 1.540 1.820 ;
        RECT  0.190 0.630 1.380 0.790 ;
        RECT  0.070 1.660 1.380 1.820 ;
    END
END AN3D1

MACRO AN3D2
    CLASS CORE ;
    FOREIGN AN3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.960 1.630 2.100 ;
        RECT  1.630 1.390 1.690 2.100 ;
        RECT  1.630 0.420 1.690 0.900 ;
        RECT  1.690 0.420 1.790 2.100 ;
        RECT  1.790 1.960 1.820 2.100 ;
        RECT  1.790 0.780 1.830 1.515 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.130 0.300 ;
        RECT  1.130 -0.300 1.350 0.340 ;
        RECT  1.350 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.700 1.510 1.800 ;
        RECT  0.430 0.700 1.350 0.840 ;
        RECT  1.070 1.680 1.350 1.800 ;
        RECT  0.850 1.680 1.070 2.100 ;
        RECT  0.290 1.680 0.850 1.800 ;
        RECT  0.210 0.420 0.430 0.840 ;
        RECT  0.070 1.680 0.290 2.100 ;
    END
END AN3D2

MACRO AN3D4
    CLASS CORE ;
    FOREIGN AN3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.650 2.830 2.030 ;
        RECT  2.500 0.490 2.830 0.870 ;
        RECT  2.830 0.490 3.250 2.030 ;
        RECT  3.250 1.650 3.410 2.030 ;
        RECT  3.250 0.490 3.410 0.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.765 0.250 1.515 ;
        RECT  0.250 0.765 1.950 0.885 ;
        RECT  1.950 0.765 2.110 1.270 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.750 1.235 ;
        RECT  0.750 1.005 0.870 1.755 ;
        RECT  0.870 1.635 1.590 1.755 ;
        RECT  1.590 1.080 1.710 1.755 ;
        RECT  1.710 1.080 1.830 1.240 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 2.090 0.300 ;
        RECT  2.090 -0.300 2.310 0.340 ;
        RECT  2.310 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 1.080 2.590 1.240 ;
        RECT  2.230 0.470 2.350 1.510 ;
        RECT  1.100 0.470 2.230 0.630 ;
        RECT  2.000 1.390 2.230 1.510 ;
        RECT  2.000 1.960 2.030 2.100 ;
        RECT  1.840 1.390 2.000 2.100 ;
        RECT  1.810 1.890 1.840 2.100 ;
        RECT  0.650 1.890 1.810 2.050 ;
        RECT  0.620 1.890 0.650 2.100 ;
        RECT  0.460 1.370 0.620 2.100 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  2.500 0.490 2.615 0.870 ;
        RECT  2.500 1.650 2.615 2.030 ;
    END
END AN3D4

MACRO AN3D8
    CLASS CORE ;
    FOREIGN AN3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.560 1.640 4.430 2.020 ;
        RECT  3.560 0.500 4.430 0.880 ;
        RECT  4.430 0.500 4.850 2.020 ;
        RECT  4.850 1.640 5.940 2.020 ;
        RECT  4.850 0.500 5.940 0.880 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.350 1.235 ;
        RECT  1.350 0.710 1.510 1.235 ;
        RECT  1.510 0.710 3.040 0.830 ;
        RECT  3.040 0.710 3.200 1.250 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.005 0.730 1.235 ;
        RECT  0.730 1.005 0.870 1.525 ;
        RECT  0.870 1.405 1.710 1.525 ;
        RECT  1.710 0.950 1.870 1.525 ;
        RECT  1.870 0.950 2.670 1.070 ;
        RECT  2.670 0.950 2.830 1.430 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.765 ;
        RECT  0.230 1.005 0.410 1.225 ;
        RECT  0.230 1.645 2.070 1.765 ;
        RECT  2.070 1.190 2.230 1.765 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 3.140 0.300 ;
        RECT  3.140 -0.300 3.360 0.340 ;
        RECT  3.360 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.440 1.100 4.215 1.260 ;
        RECT  3.320 0.470 3.440 1.745 ;
        RECT  2.370 0.470 3.320 0.590 ;
        RECT  3.060 1.625 3.320 1.745 ;
        RECT  2.840 1.625 3.060 2.045 ;
        RECT  0.070 1.885 2.840 2.045 ;
        RECT  2.150 0.430 2.370 0.590 ;
        RECT  0.290 0.470 2.150 0.590 ;
        RECT  0.070 0.470 0.290 0.885 ;
        LAYER M1 ;
        RECT  3.560 0.500 4.215 0.880 ;
        RECT  3.560 1.640 4.215 2.020 ;
        RECT  5.065 0.500 5.940 0.880 ;
        RECT  5.065 1.640 5.940 2.020 ;
    END
END AN3D8

MACRO AN4D0
    CLASS CORE ;
    FOREIGN AN4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.520 2.150 1.810 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.990 1.520 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.990 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.990 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.990 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.520 0.300 ;
        RECT  1.520 -0.300 1.740 0.340 ;
        RECT  1.740 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.795 2.820 ;
        RECT  0.795 2.180 1.015 2.820 ;
        RECT  1.015 2.220 1.550 2.820 ;
        RECT  1.550 2.180 1.770 2.820 ;
        RECT  1.770 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.710 0.570 1.870 1.795 ;
        RECT  0.430 1.635 1.710 1.795 ;
        RECT  0.190 0.570 1.710 0.730 ;
    END
END AN4D0

MACRO AN4D1
    CLASS CORE ;
    FOREIGN AN4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  1.990 0.420 2.150 2.100 ;
        RECT  2.150 1.960 2.180 2.100 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.990 1.520 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.990 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.990 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.990 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.510 0.300 ;
        RECT  1.510 -0.300 1.730 0.340 ;
        RECT  1.730 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.795 2.820 ;
        RECT  0.795 2.180 1.015 2.820 ;
        RECT  1.015 2.220 1.550 2.820 ;
        RECT  1.550 2.180 1.770 2.820 ;
        RECT  1.770 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.570 1.850 1.795 ;
        RECT  0.190 0.570 1.690 0.730 ;
        RECT  0.430 1.635 1.690 1.795 ;
    END
END AN4D1

MACRO AN4D2
    CLASS CORE ;
    FOREIGN AN4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.950 1.390 2.010 2.100 ;
        RECT  1.950 0.420 2.010 0.900 ;
        RECT  2.010 0.420 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.780 2.150 1.515 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.520 0.300 ;
        RECT  1.520 -0.300 1.740 0.340 ;
        RECT  1.740 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.820 1.080 1.840 1.240 ;
        RECT  1.680 0.690 1.820 1.800 ;
        RECT  0.440 0.690 1.680 0.850 ;
        RECT  1.390 1.640 1.680 1.800 ;
        RECT  1.170 1.640 1.390 2.060 ;
        RECT  0.690 1.640 1.170 1.800 ;
        RECT  0.470 1.640 0.690 2.060 ;
        RECT  0.220 0.430 0.440 0.850 ;
    END
END AN4D2

MACRO AN4D4
    CLASS CORE ;
    FOREIGN AN4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.250 1.640 3.790 2.020 ;
        RECT  3.250 0.500 3.790 0.880 ;
        RECT  3.790 0.500 4.210 2.020 ;
        RECT  4.210 1.640 4.270 2.020 ;
        RECT  4.210 0.500 4.270 0.880 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 0.765 0.490 1.270 ;
        RECT  0.490 0.765 2.650 0.885 ;
        RECT  2.650 0.765 2.810 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.080 0.730 1.240 ;
        RECT  0.730 1.080 0.850 1.755 ;
        RECT  0.850 1.635 2.310 1.755 ;
        RECT  2.310 1.005 2.470 1.755 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.030 1.150 1.515 ;
        RECT  1.150 1.395 1.990 1.515 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.650 0.300 ;
        RECT  3.650 -0.300 3.870 0.340 ;
        RECT  3.870 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.650 2.820 ;
        RECT  3.650 2.180 3.870 2.820 ;
        RECT  3.870 2.220 4.450 2.820 ;
        RECT  4.450 2.180 4.670 2.820 ;
        RECT  4.670 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.090 1.080 3.360 1.240 ;
        RECT  2.970 0.470 3.090 2.050 ;
        RECT  1.470 0.470 2.970 0.630 ;
        RECT  0.640 1.890 2.970 2.050 ;
        RECT  0.610 1.890 0.640 2.100 ;
        RECT  0.450 1.390 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  3.250 0.500 3.575 0.880 ;
        RECT  3.250 1.640 3.575 2.020 ;
    END
END AN4D4

MACRO AN4D8
    CLASS CORE ;
    FOREIGN AN4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.900 1.640 6.030 2.020 ;
        RECT  4.870 0.500 6.030 0.880 ;
        RECT  6.030 0.500 6.450 2.020 ;
        RECT  6.450 1.640 7.260 2.020 ;
        RECT  6.450 0.500 7.260 0.880 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 4.070 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.230 2.820 ;
        RECT  2.230 2.180 2.450 2.820 ;
        RECT  2.450 2.220 3.030 2.820 ;
        RECT  3.030 2.180 3.250 2.820 ;
        RECT  3.250 2.220 4.510 2.820 ;
        RECT  4.510 2.180 4.730 2.820 ;
        RECT  4.730 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.570 0.750 3.350 0.870 ;
        RECT  2.350 0.450 2.570 0.870 ;
        RECT  4.180 0.470 4.400 0.850 ;
        RECT  3.710 0.470 4.180 0.630 ;
        RECT  3.490 0.470 3.710 0.850 ;
        RECT  4.555 1.080 5.490 1.240 ;
        RECT  4.435 1.080 4.555 1.500 ;
        RECT  4.310 1.380 4.435 1.500 ;
        RECT  4.310 1.930 4.340 2.090 ;
        RECT  4.150 1.380 4.310 2.090 ;
        RECT  3.620 1.380 4.150 1.500 ;
        RECT  4.120 1.930 4.150 2.090 ;
        RECT  3.620 1.930 3.650 2.090 ;
        RECT  3.460 1.380 3.620 2.090 ;
        RECT  2.820 1.380 3.460 1.500 ;
        RECT  3.430 1.930 3.460 2.090 ;
        RECT  2.820 1.930 2.850 2.090 ;
        RECT  2.660 1.380 2.820 2.090 ;
        RECT  2.020 1.380 2.660 1.500 ;
        RECT  2.630 1.930 2.660 2.090 ;
        RECT  2.020 1.930 2.050 2.090 ;
        RECT  1.860 1.380 2.020 2.090 ;
        RECT  1.330 1.380 1.860 1.500 ;
        RECT  1.830 1.930 1.860 2.090 ;
        RECT  1.330 1.930 1.360 2.090 ;
        RECT  1.170 1.380 1.330 2.090 ;
        RECT  1.050 1.380 1.170 1.500 ;
        RECT  1.140 1.930 1.170 2.090 ;
        RECT  0.910 0.750 1.050 1.500 ;
        RECT  0.290 0.750 0.910 0.870 ;
        RECT  0.640 1.380 0.910 1.500 ;
        RECT  0.640 1.930 0.670 2.090 ;
        RECT  0.480 1.380 0.640 2.090 ;
        RECT  0.450 1.930 0.480 2.090 ;
        RECT  2.710 0.470 3.490 0.630 ;
        RECT  1.570 0.750 2.350 0.870 ;
        RECT  0.070 0.470 0.290 0.870 ;
        RECT  0.430 0.470 2.210 0.630 ;
        LAYER M1 ;
        RECT  4.870 0.500 5.815 0.880 ;
        RECT  4.900 1.640 5.815 2.020 ;
        RECT  6.665 0.500 7.260 0.880 ;
        RECT  6.665 1.640 7.260 2.020 ;
    END
END AN4D8

MACRO ANTENNA
    CLASS CORE ;
    FOREIGN ANTENNA 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.795 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
END ANTENNA

MACRO AO211D0
    CLASS CORE ;
    FOREIGN AO211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.660 2.150 1.710 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.080 0.720 1.240 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.080 1.050 1.240 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.720 0.300 ;
        RECT  0.720 -0.300 0.940 0.340 ;
        RECT  0.940 -0.300 1.670 0.300 ;
        RECT  1.670 -0.300 1.890 0.340 ;
        RECT  1.890 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.670 2.820 ;
        RECT  1.670 2.180 1.890 2.820 ;
        RECT  1.890 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 0.710 1.850 1.795 ;
        RECT  0.350 0.710 1.690 0.870 ;
        RECT  0.970 1.635 1.690 1.795 ;
    END
END AO211D0

MACRO AO211D1
    CLASS CORE ;
    FOREIGN AO211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  1.990 0.420 2.150 2.100 ;
        RECT  2.150 1.960 2.180 2.100 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.280 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.790 0.300 ;
        RECT  0.790 -0.300 1.010 0.340 ;
        RECT  1.010 -0.300 1.570 0.300 ;
        RECT  1.570 -0.300 1.790 0.340 ;
        RECT  1.790 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.550 2.820 ;
        RECT  1.550 2.180 1.770 2.820 ;
        RECT  1.770 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.370 0.750 1.180 0.870 ;
        RECT  1.180 0.450 1.400 0.870 ;
        RECT  0.440 1.635 1.700 1.795 ;
        RECT  1.400 0.750 1.700 0.870 ;
        RECT  1.700 0.750 1.860 1.795 ;
        RECT  0.100 1.370 0.260 2.095 ;
        RECT  0.260 1.915 0.290 2.095 ;
        RECT  0.290 1.915 0.860 2.035 ;
        RECT  0.860 1.915 1.100 2.075 ;
        RECT  0.070 1.960 0.100 2.095 ;
        RECT  0.150 0.450 0.370 0.870 ;
    END
END AO211D1

MACRO AO211D2
    CLASS CORE ;
    FOREIGN AO211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.950 1.390 2.010 2.100 ;
        RECT  1.950 0.420 2.010 0.900 ;
        RECT  2.010 0.420 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.780 2.150 1.515 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.710 0.300 ;
        RECT  0.710 -0.300 0.930 0.340 ;
        RECT  0.930 -0.300 1.520 0.300 ;
        RECT  1.520 -0.300 1.740 0.340 ;
        RECT  1.740 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.530 2.820 ;
        RECT  1.530 2.180 1.750 2.820 ;
        RECT  1.750 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 1.915 0.860 2.035 ;
        RECT  0.860 1.915 1.100 2.075 ;
        RECT  0.260 1.915 0.290 2.095 ;
        RECT  0.100 1.370 0.260 2.095 ;
        RECT  1.830 1.070 1.850 1.240 ;
        RECT  1.690 0.750 1.830 1.795 ;
        RECT  1.330 0.750 1.690 0.870 ;
        RECT  0.440 1.635 1.690 1.795 ;
        RECT  1.110 0.450 1.330 0.870 ;
        RECT  0.280 0.750 1.110 0.870 ;
        RECT  0.060 0.450 0.280 0.870 ;
        RECT  0.070 1.960 0.100 2.095 ;
    END
END AO211D2

MACRO AO211D4
    CLASS CORE ;
    FOREIGN AO211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.650 3.790 2.030 ;
        RECT  3.610 0.490 3.790 0.870 ;
        RECT  3.790 0.490 4.210 2.030 ;
        RECT  4.210 1.650 4.610 2.030 ;
        RECT  4.210 0.490 4.610 0.870 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.765 0.250 1.515 ;
        RECT  0.250 0.765 1.230 0.885 ;
        RECT  1.230 0.765 1.390 1.270 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.660 0.765 1.820 1.270 ;
        RECT  1.820 0.765 2.650 0.885 ;
        RECT  2.650 0.765 2.770 1.240 ;
        RECT  2.770 1.005 3.110 1.240 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.240 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.330 ;
        RECT  2.990 -0.300 3.210 0.300 ;
        RECT  3.210 -0.300 3.430 0.340 ;
        RECT  3.430 -0.300 4.000 0.300 ;
        RECT  4.000 -0.300 4.220 0.330 ;
        RECT  4.220 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.330 ;
        RECT  5.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.700 2.820 ;
        RECT  0.700 2.180 0.920 2.820 ;
        RECT  0.920 2.220 3.220 2.820 ;
        RECT  3.220 2.180 3.440 2.820 ;
        RECT  3.440 2.220 4.000 2.820 ;
        RECT  4.000 2.180 4.220 2.820 ;
        RECT  4.220 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.870 1.680 3.090 2.100 ;
        RECT  2.330 1.890 2.870 2.050 ;
        RECT  2.110 1.680 2.330 2.100 ;
        RECT  1.570 1.890 2.110 2.050 ;
        RECT  1.540 1.890 1.570 2.100 ;
        RECT  1.380 1.390 1.540 2.100 ;
        RECT  1.350 1.890 1.380 2.100 ;
        RECT  0.280 1.890 1.350 2.050 ;
        RECT  3.240 0.470 3.400 1.560 ;
        RECT  0.400 0.470 3.240 0.630 ;
        RECT  1.730 1.400 3.240 1.560 ;
        RECT  0.060 1.635 0.280 2.050 ;
        LAYER M1 ;
        RECT  4.425 0.490 4.610 0.870 ;
        RECT  4.425 1.650 4.610 2.030 ;
    END
END AO211D4

MACRO AO21D0
    CLASS CORE ;
    FOREIGN AO21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.420 1.830 1.930 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.285 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.220 0.300 ;
        RECT  1.220 -0.300 1.440 0.340 ;
        RECT  1.440 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.230 2.820 ;
        RECT  1.230 2.180 1.450 2.820 ;
        RECT  1.450 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 1.670 1.020 2.050 ;
        RECT  0.260 1.930 0.860 2.050 ;
        RECT  1.360 0.470 1.520 1.270 ;
        RECT  1.020 0.470 1.360 0.590 ;
        RECT  0.800 0.430 1.020 0.590 ;
        RECT  0.570 0.470 0.800 0.590 ;
        RECT  0.100 1.670 0.260 2.050 ;
        RECT  0.450 0.470 0.570 1.810 ;
        RECT  0.570 1.660 0.690 1.810 ;
    END
END AO21D0

MACRO AO21D1
    CLASS CORE ;
    FOREIGN AO21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.670 0.420 1.830 2.100 ;
        RECT  1.830 1.960 1.860 2.100 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.230 0.300 ;
        RECT  1.230 -0.300 1.450 0.340 ;
        RECT  1.450 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.240 2.820 ;
        RECT  1.240 2.180 1.460 2.820 ;
        RECT  1.460 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  0.830 1.635 1.050 2.075 ;
        RECT  1.390 0.745 1.550 1.290 ;
        RECT  1.010 0.745 1.390 0.885 ;
        RECT  0.790 0.470 1.010 0.885 ;
        RECT  0.570 0.745 0.790 0.885 ;
        RECT  0.570 1.630 0.670 1.790 ;
        RECT  0.450 0.745 0.570 1.790 ;
        RECT  0.070 1.635 0.290 2.075 ;
    END
END AO21D1

MACRO AO21D2
    CLASS CORE ;
    FOREIGN AO21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.960 1.630 2.100 ;
        RECT  1.630 1.390 1.690 2.100 ;
        RECT  1.630 0.420 1.690 0.900 ;
        RECT  1.690 0.420 1.790 2.100 ;
        RECT  1.790 1.960 1.820 2.100 ;
        RECT  1.790 0.780 1.830 1.515 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.210 0.300 ;
        RECT  1.210 -0.300 1.430 0.340 ;
        RECT  1.430 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 1.635 1.050 2.075 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  1.510 1.050 1.530 1.290 ;
        RECT  1.370 0.745 1.510 1.290 ;
        RECT  1.010 0.745 1.370 0.885 ;
        RECT  0.790 0.470 1.010 0.885 ;
        RECT  0.570 0.745 0.790 0.885 ;
        RECT  0.570 1.630 0.670 1.790 ;
        RECT  0.070 1.635 0.290 2.075 ;
        RECT  0.450 0.745 0.570 1.790 ;
    END
END AO21D2

MACRO AO21D4
    CLASS CORE ;
    FOREIGN AO21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.650 3.150 2.030 ;
        RECT  2.630 0.490 3.150 0.870 ;
        RECT  3.150 0.490 3.570 2.030 ;
        RECT  3.570 1.650 3.640 2.030 ;
        RECT  3.570 0.490 3.640 0.870 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        RECT  0.230 1.005 0.370 1.240 ;
        RECT  0.370 0.765 0.490 1.240 ;
        RECT  0.490 0.765 2.100 0.885 ;
        RECT  2.100 0.765 2.260 1.290 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.030 0.840 1.490 ;
        RECT  0.840 1.370 1.690 1.490 ;
        RECT  1.690 1.005 1.830 1.490 ;
        RECT  1.830 1.050 1.900 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 2.240 0.300 ;
        RECT  2.240 -0.300 2.460 0.340 ;
        RECT  2.460 -0.300 3.020 0.300 ;
        RECT  3.020 -0.300 3.240 0.340 ;
        RECT  3.240 -0.300 3.810 0.300 ;
        RECT  3.810 -0.300 4.030 0.340 ;
        RECT  4.030 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 3.810 2.820 ;
        RECT  3.810 2.180 4.030 2.820 ;
        RECT  4.030 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.640 1.890 2.180 2.050 ;
        RECT  2.510 1.080 2.740 1.240 ;
        RECT  2.390 0.470 2.510 1.770 ;
        RECT  0.500 0.470 2.390 0.630 ;
        RECT  0.780 1.610 2.390 1.770 ;
        RECT  0.420 1.630 0.640 2.050 ;
        LAYER M1 ;
        RECT  2.630 0.490 2.935 0.870 ;
        RECT  2.630 1.650 2.935 2.030 ;
    END
END AO21D4

MACRO AO221D0
    CLASS CORE ;
    FOREIGN AO221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.420 2.470 1.860 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.255 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.720 0.240 1.515 ;
        RECT  0.240 0.720 1.030 0.860 ;
        RECT  1.030 0.720 1.250 0.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.520 1.260 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.980 0.570 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.100 0.340 ;
        RECT  1.100 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.950 2.820 ;
        RECT  1.950 2.180 2.170 2.820 ;
        RECT  2.170 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.790 1.650 1.220 1.810 ;
        RECT  1.220 1.380 1.340 1.810 ;
        RECT  0.440 0.470 1.540 0.600 ;
        RECT  1.540 0.440 1.760 0.600 ;
        RECT  1.340 1.380 2.050 1.500 ;
        RECT  1.760 0.470 2.050 0.600 ;
        RECT  2.050 0.470 2.190 1.500 ;
        RECT  0.500 1.650 0.620 2.050 ;
        RECT  0.620 1.930 1.580 2.050 ;
        RECT  1.580 1.620 1.740 2.050 ;
        RECT  0.070 1.650 0.500 1.810 ;
        RECT  0.200 0.440 0.440 0.600 ;
    END
END AO221D0

MACRO AO221D1
    CLASS CORE ;
    FOREIGN AO221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 1.420 2.650 2.100 ;
        RECT  2.630 0.420 2.650 0.870 ;
        RECT  2.650 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.190 1.270 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.130 0.300 ;
        RECT  1.130 -0.300 1.350 0.340 ;
        RECT  1.350 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 0.730 1.790 0.850 ;
        RECT  1.790 0.430 2.010 0.850 ;
        RECT  2.010 0.730 2.380 0.850 ;
        RECT  2.380 0.730 2.500 1.290 ;
        RECT  2.500 1.050 2.530 1.290 ;
        RECT  1.340 1.910 1.880 2.050 ;
        RECT  1.880 1.650 2.100 2.070 ;
        RECT  0.290 1.930 0.860 2.050 ;
        RECT  0.860 1.450 1.000 2.050 ;
        RECT  1.000 1.450 1.020 1.790 ;
        RECT  1.020 1.635 1.740 1.790 ;
        RECT  0.760 0.430 0.980 0.850 ;
        RECT  0.570 0.730 0.760 0.850 ;
        RECT  0.570 1.400 0.670 1.810 ;
        RECT  1.120 1.910 1.340 2.070 ;
        RECT  0.070 1.650 0.290 2.070 ;
        RECT  0.450 0.730 0.570 1.810 ;
    END
END AO221D1

MACRO AO221D2
    CLASS CORE ;
    FOREIGN AO221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.960 2.590 2.100 ;
        RECT  2.590 1.390 2.650 2.100 ;
        RECT  2.590 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.750 2.100 ;
        RECT  2.750 1.960 2.780 2.100 ;
        RECT  2.750 0.780 2.790 1.515 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.190 1.270 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.005 1.510 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.130 0.300 ;
        RECT  1.130 -0.300 1.350 0.340 ;
        RECT  1.350 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.020 1.635 1.730 1.790 ;
        RECT  0.980 1.450 1.020 1.790 ;
        RECT  0.860 1.450 0.980 2.050 ;
        RECT  0.290 1.930 0.860 2.050 ;
        RECT  1.870 1.650 2.090 2.070 ;
        RECT  1.330 1.910 1.870 2.050 ;
        RECT  2.470 1.050 2.530 1.270 ;
        RECT  2.350 0.760 2.470 1.270 ;
        RECT  2.010 0.760 2.350 0.880 ;
        RECT  1.790 0.430 2.010 0.880 ;
        RECT  0.980 0.760 1.790 0.880 ;
        RECT  0.760 0.430 0.980 0.880 ;
        RECT  0.570 0.760 0.760 0.880 ;
        RECT  0.570 1.400 0.670 1.810 ;
        RECT  0.450 0.760 0.570 1.810 ;
        RECT  1.110 1.910 1.330 2.070 ;
        RECT  0.070 1.650 0.290 2.070 ;
    END
END AO221D2

MACRO AO221D4
    CLASS CORE ;
    FOREIGN AO221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.800 1.650 5.070 2.030 ;
        RECT  4.800 0.490 5.070 0.870 ;
        RECT  5.070 0.490 5.490 2.030 ;
        RECT  5.490 1.650 5.840 2.030 ;
        RECT  5.490 0.490 5.840 0.870 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.100 1.240 ;
        RECT  1.100 1.005 1.220 1.480 ;
        RECT  1.220 1.360 2.110 1.480 ;
        RECT  2.110 1.030 2.270 1.480 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.990 1.235 ;
        RECT  2.990 1.005 3.110 1.475 ;
        RECT  3.110 1.355 3.900 1.475 ;
        RECT  3.900 1.030 4.060 1.475 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.570 0.300 ;
        RECT  1.570 -0.300 1.790 0.340 ;
        RECT  1.790 -0.300 3.350 0.300 ;
        RECT  3.350 -0.300 3.570 0.340 ;
        RECT  3.570 -0.300 4.410 0.300 ;
        RECT  4.410 -0.300 4.630 0.340 ;
        RECT  4.630 -0.300 5.210 0.300 ;
        RECT  5.210 -0.300 5.430 0.340 ;
        RECT  5.430 -0.300 6.030 0.300 ;
        RECT  6.030 -0.300 6.250 0.340 ;
        RECT  6.250 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.210 2.820 ;
        RECT  5.210 2.180 5.430 2.820 ;
        RECT  5.430 2.220 6.030 2.820 ;
        RECT  6.030 2.180 6.250 2.820 ;
        RECT  6.250 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 1.890 2.510 2.050 ;
        RECT  0.960 1.890 0.990 2.100 ;
        RECT  0.800 1.370 0.960 2.100 ;
        RECT  0.770 1.890 0.800 2.100 ;
        RECT  0.250 1.890 0.770 2.050 ;
        RECT  4.520 0.770 4.680 1.510 ;
        RECT  4.240 0.770 4.520 0.890 ;
        RECT  4.340 1.390 4.520 1.510 ;
        RECT  4.340 1.960 4.370 2.100 ;
        RECT  4.180 1.390 4.340 2.100 ;
        RECT  4.020 0.470 4.240 0.890 ;
        RECT  4.150 1.890 4.180 2.100 ;
        RECT  2.630 1.890 4.150 2.050 ;
        RECT  2.910 0.470 4.020 0.630 ;
        RECT  2.690 0.470 2.910 0.885 ;
        RECT  2.460 0.470 2.690 0.630 ;
        RECT  2.240 0.470 2.460 0.890 ;
        RECT  1.130 0.470 2.240 0.630 ;
        RECT  0.910 0.470 1.130 0.885 ;
        RECT  0.300 0.470 0.910 0.630 ;
        RECT  1.130 1.610 4.010 1.770 ;
        RECT  0.090 1.550 0.250 2.050 ;
        RECT  0.080 0.470 0.300 0.890 ;
        LAYER M1 ;
        RECT  4.800 0.490 4.855 0.870 ;
        RECT  4.800 1.650 4.855 2.030 ;
        RECT  5.700 0.490 5.840 0.870 ;
        RECT  5.705 1.650 5.840 2.030 ;
    END
END AO221D4

MACRO AO222D0
    CLASS CORE ;
    FOREIGN AO222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 0.660 3.110 1.710 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.255 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.720 0.240 1.515 ;
        RECT  0.240 0.720 1.030 0.840 ;
        RECT  1.030 0.720 1.250 0.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.530 1.255 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.960 0.570 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.870 0.300 ;
        RECT  0.870 -0.300 1.090 0.340 ;
        RECT  1.090 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.910 2.820 ;
        RECT  1.910 2.180 2.130 2.820 ;
        RECT  2.130 2.220 2.630 2.820 ;
        RECT  2.630 2.180 2.850 2.820 ;
        RECT  2.850 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.670 1.650 2.510 1.810 ;
        RECT  1.550 1.650 1.670 2.050 ;
        RECT  0.620 1.930 1.550 2.050 ;
        RECT  0.500 1.650 0.620 2.050 ;
        RECT  2.650 0.470 2.810 1.530 ;
        RECT  1.760 0.470 2.650 0.590 ;
        RECT  1.340 1.410 2.650 1.530 ;
        RECT  1.540 0.430 1.760 0.590 ;
        RECT  0.430 0.470 1.540 0.590 ;
        RECT  1.220 1.410 1.340 1.810 ;
        RECT  0.790 1.650 1.220 1.810 ;
        RECT  0.070 1.650 0.500 1.810 ;
        RECT  0.190 0.430 0.430 0.590 ;
    END
END AO222D0

MACRO AO222D1
    CLASS CORE ;
    FOREIGN AO222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.960 2.950 2.100 ;
        RECT  2.950 1.390 2.990 2.100 ;
        RECT  2.940 0.420 2.990 0.900 ;
        RECT  2.990 0.420 3.110 2.100 ;
        RECT  3.110 1.960 3.140 2.100 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.550 1.270 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 1.490 0.300 ;
        RECT  1.490 -0.300 1.710 0.340 ;
        RECT  1.710 -0.300 2.510 0.300 ;
        RECT  2.510 -0.300 2.730 0.340 ;
        RECT  2.730 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.700 0.725 2.820 1.290 ;
        RECT  2.820 1.050 2.870 1.290 ;
        RECT  2.230 1.635 2.450 2.070 ;
        RECT  0.290 1.910 0.830 2.050 ;
        RECT  0.830 1.650 1.050 2.070 ;
        RECT  1.050 1.910 1.590 2.050 ;
        RECT  1.590 1.910 1.830 2.070 ;
        RECT  2.070 0.725 2.700 0.855 ;
        RECT  1.850 0.435 2.070 0.855 ;
        RECT  1.060 0.725 1.850 0.855 ;
        RECT  0.840 0.435 1.060 0.855 ;
        RECT  0.220 0.725 0.840 0.855 ;
        RECT  0.220 1.635 0.690 1.790 ;
        RECT  0.100 0.725 0.220 1.790 ;
        RECT  1.190 1.635 2.230 1.790 ;
        RECT  0.070 1.910 0.290 2.070 ;
    END
END AO222D1

MACRO AO222D2
    CLASS CORE ;
    FOREIGN AO222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.090 1.960 3.120 2.100 ;
        RECT  3.000 0.420 3.170 0.900 ;
        RECT  3.120 1.390 3.280 2.100 ;
        RECT  3.280 1.390 3.290 1.515 ;
        RECT  3.170 0.780 3.290 0.900 ;
        RECT  3.280 1.960 3.310 2.100 ;
        RECT  3.290 0.780 3.430 1.515 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.630 1.240 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 1.490 0.300 ;
        RECT  1.490 -0.300 1.710 0.340 ;
        RECT  1.710 -0.300 2.570 0.300 ;
        RECT  2.570 -0.300 2.790 0.340 ;
        RECT  2.790 -0.300 3.380 0.300 ;
        RECT  3.380 -0.300 3.600 0.340 ;
        RECT  3.600 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.690 2.820 ;
        RECT  2.690 2.180 2.910 2.820 ;
        RECT  2.910 2.220 3.490 2.820 ;
        RECT  3.490 2.180 3.710 2.820 ;
        RECT  3.710 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.590 1.910 1.830 2.070 ;
        RECT  1.050 1.910 1.590 2.050 ;
        RECT  0.830 1.650 1.050 2.070 ;
        RECT  0.290 1.910 0.830 2.050 ;
        RECT  2.290 1.635 2.510 2.070 ;
        RECT  2.880 1.080 3.060 1.240 ;
        RECT  2.760 0.725 2.880 1.240 ;
        RECT  2.130 0.725 2.760 0.855 ;
        RECT  1.910 0.435 2.130 0.855 ;
        RECT  1.060 0.725 1.910 0.855 ;
        RECT  0.840 0.435 1.060 0.855 ;
        RECT  0.220 0.725 0.840 0.855 ;
        RECT  0.220 1.635 0.690 1.790 ;
        RECT  1.190 1.635 2.290 1.790 ;
        RECT  0.100 0.725 0.220 1.790 ;
        RECT  0.070 1.910 0.290 2.070 ;
    END
END AO222D2

MACRO AO222D4
    CLASS CORE ;
    FOREIGN AO222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.630 1.650 6.030 2.030 ;
        RECT  5.630 0.490 6.030 0.870 ;
        RECT  6.030 0.490 6.450 2.030 ;
        RECT  6.450 1.650 6.580 2.030 ;
        RECT  6.450 0.490 6.580 0.870 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.395 1.380 1.515 ;
        RECT  1.380 1.030 1.540 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.515 ;
        RECT  2.150 1.395 2.910 1.515 ;
        RECT  2.910 1.030 3.070 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.515 ;
        RECT  3.750 1.395 4.700 1.515 ;
        RECT  4.700 1.030 4.860 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.210 0.300 ;
        RECT  0.210 -0.300 0.430 0.340 ;
        RECT  0.430 -0.300 1.530 0.300 ;
        RECT  1.530 -0.300 1.750 0.340 ;
        RECT  1.750 -0.300 2.980 0.300 ;
        RECT  2.980 -0.300 3.200 0.340 ;
        RECT  3.200 -0.300 4.150 0.300 ;
        RECT  4.150 -0.300 4.370 0.340 ;
        RECT  4.370 -0.300 5.220 0.300 ;
        RECT  5.220 -0.300 5.440 0.340 ;
        RECT  5.440 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.790 1.635 3.310 1.795 ;
        RECT  1.570 1.635 1.790 2.055 ;
        RECT  1.090 1.635 1.570 1.795 ;
        RECT  0.870 1.635 1.090 2.055 ;
        RECT  0.290 1.635 0.870 1.795 ;
        RECT  4.570 1.915 4.810 2.075 ;
        RECT  4.030 1.915 4.570 2.035 ;
        RECT  3.810 1.915 4.030 2.075 ;
        RECT  2.930 1.915 3.810 2.035 ;
        RECT  2.710 1.915 2.930 2.075 ;
        RECT  2.170 1.915 2.710 2.035 ;
        RECT  5.480 1.080 5.740 1.240 ;
        RECT  5.360 0.765 5.480 1.795 ;
        RECT  5.040 0.765 5.360 0.885 ;
        RECT  5.170 1.635 5.360 1.795 ;
        RECT  4.950 1.635 5.170 2.055 ;
        RECT  4.820 0.470 5.040 0.885 ;
        RECT  3.430 1.635 4.950 1.795 ;
        RECT  3.710 0.765 4.820 0.885 ;
        RECT  3.490 0.470 3.710 0.885 ;
        RECT  2.420 0.765 3.490 0.885 ;
        RECT  2.200 0.470 2.420 0.885 ;
        RECT  1.090 0.765 2.200 0.885 ;
        RECT  1.930 1.915 2.170 2.075 ;
        RECT  0.070 1.635 0.290 2.055 ;
        RECT  0.870 0.470 1.090 0.885 ;
        LAYER M1 ;
        RECT  5.630 0.490 5.815 0.870 ;
        RECT  5.630 1.650 5.815 2.030 ;
    END
END AO222D4

MACRO AO22D0
    CLASS CORE ;
    FOREIGN AO22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.440 2.150 2.040 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 0.725 0.700 1.150 ;
        RECT  0.700 0.725 1.370 0.845 ;
        RECT  1.370 0.725 1.510 1.235 ;
        RECT  1.510 0.940 1.600 1.160 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.190 1.250 1.410 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.285 0.870 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.535 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.460 0.300 ;
        RECT  1.460 -0.300 1.680 0.340 ;
        RECT  1.680 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.220 1.930 1.460 2.090 ;
        RECT  0.660 1.930 1.220 2.050 ;
        RECT  1.720 0.485 1.870 1.810 ;
        RECT  0.930 0.485 1.720 0.605 ;
        RECT  0.810 1.650 1.720 1.810 ;
        RECT  0.420 1.930 0.660 2.090 ;
        RECT  0.690 0.445 0.930 0.605 ;
    END
END AO22D0

MACRO AO22D1
    CLASS CORE ;
    FOREIGN AO22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.960 2.310 2.100 ;
        RECT  2.310 0.420 2.470 2.100 ;
        RECT  2.470 1.960 2.500 2.100 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.800 0.300 ;
        RECT  0.800 -0.300 1.020 0.340 ;
        RECT  1.020 -0.300 1.870 0.300 ;
        RECT  1.870 -0.300 2.090 0.340 ;
        RECT  2.090 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.890 2.820 ;
        RECT  1.890 2.180 2.110 2.820 ;
        RECT  2.110 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.545 1.910 1.780 2.070 ;
        RECT  1.000 1.910 1.545 2.050 ;
        RECT  0.780 1.635 1.000 2.050 ;
        RECT  0.280 1.910 0.780 2.050 ;
        RECT  1.980 0.765 2.140 1.790 ;
        RECT  1.690 0.765 1.980 0.885 ;
        RECT  1.140 1.635 1.980 1.790 ;
        RECT  1.470 0.470 1.690 0.885 ;
        RECT  0.360 0.765 1.470 0.885 ;
        RECT  0.140 0.470 0.360 0.885 ;
        RECT  0.060 1.635 0.280 2.050 ;
    END
END AO22D1

MACRO AO22D2
    CLASS CORE ;
    FOREIGN AO22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.960 2.270 2.100 ;
        RECT  2.270 1.390 2.330 2.100 ;
        RECT  2.270 0.420 2.330 0.900 ;
        RECT  2.330 0.420 2.430 2.100 ;
        RECT  2.430 1.960 2.460 2.100 ;
        RECT  2.430 0.780 2.470 1.515 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.800 0.300 ;
        RECT  0.800 -0.300 1.020 0.340 ;
        RECT  1.020 -0.300 1.850 0.300 ;
        RECT  1.850 -0.300 2.070 0.340 ;
        RECT  2.070 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.545 1.910 1.780 2.070 ;
        RECT  1.000 1.910 1.545 2.050 ;
        RECT  0.780 1.635 1.000 2.050 ;
        RECT  0.280 1.910 0.780 2.050 ;
        RECT  1.990 0.765 2.150 1.790 ;
        RECT  1.690 0.765 1.990 0.885 ;
        RECT  1.140 1.635 1.990 1.790 ;
        RECT  1.470 0.470 1.690 0.885 ;
        RECT  0.360 0.765 1.470 0.885 ;
        RECT  0.140 0.470 0.360 0.885 ;
        RECT  0.060 1.635 0.280 2.050 ;
    END
END AO22D2

MACRO AO22D4
    CLASS CORE ;
    FOREIGN AO22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.650 4.110 2.030 ;
        RECT  3.750 0.490 4.110 0.870 ;
        RECT  4.110 0.490 4.530 2.030 ;
        RECT  4.530 1.650 4.680 2.030 ;
        RECT  4.530 0.490 4.680 0.870 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.475 ;
        RECT  2.150 1.355 2.910 1.475 ;
        RECT  2.910 1.030 3.070 1.475 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        RECT  0.570 1.395 1.390 1.515 ;
        RECT  1.390 1.030 1.550 1.515 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.220 0.300 ;
        RECT  0.220 -0.300 0.440 0.340 ;
        RECT  0.440 -0.300 1.600 0.300 ;
        RECT  1.600 -0.300 1.820 0.340 ;
        RECT  1.820 -0.300 2.970 0.300 ;
        RECT  2.970 -0.300 3.190 0.340 ;
        RECT  3.190 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.790 1.890 3.330 2.050 ;
        RECT  1.570 1.635 1.790 2.050 ;
        RECT  1.100 1.930 1.570 2.050 ;
        RECT  0.880 1.635 1.100 2.050 ;
        RECT  0.280 1.930 0.880 2.050 ;
        RECT  0.250 1.930 0.280 2.100 ;
        RECT  0.090 1.370 0.250 2.100 ;
        RECT  3.435 0.765 3.595 1.770 ;
        RECT  2.550 0.765 3.435 0.885 ;
        RECT  1.930 1.610 3.435 1.770 ;
        RECT  2.330 0.470 2.550 0.885 ;
        RECT  1.100 0.765 2.330 0.885 ;
        RECT  0.880 0.470 1.100 0.885 ;
        RECT  0.060 1.960 0.090 2.100 ;
        LAYER M1 ;
        RECT  3.750 0.490 3.895 0.870 ;
        RECT  3.750 1.650 3.895 2.030 ;
    END
END AO22D4

MACRO AO31D0
    CLASS CORE ;
    FOREIGN AO31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.480 2.150 1.980 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 0.990 1.050 1.230 ;
        RECT  1.050 0.990 1.190 1.515 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 0.990 1.520 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.490 0.300 ;
        RECT  1.490 -0.300 1.710 0.340 ;
        RECT  1.710 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 1.880 1.450 2.050 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  1.715 0.530 1.870 1.760 ;
        RECT  1.050 0.530 1.715 0.690 ;
        RECT  1.050 1.640 1.715 1.760 ;
        RECT  0.830 1.640 1.050 1.810 ;
        RECT  0.260 1.640 0.830 1.760 ;
        RECT  0.430 1.880 0.670 2.050 ;
        RECT  0.100 1.640 0.260 1.980 ;
    END
END AO31D0

MACRO AO31D1
    CLASS CORE ;
    FOREIGN AO31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  1.990 0.420 2.150 2.100 ;
        RECT  2.150 1.960 2.180 2.100 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.540 0.300 ;
        RECT  1.540 -0.300 1.760 0.340 ;
        RECT  1.760 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 1.915 1.450 2.075 ;
        RECT  0.670 1.915 1.210 2.050 ;
        RECT  1.710 0.765 1.870 1.795 ;
        RECT  1.340 0.765 1.710 0.885 ;
        RECT  0.260 1.635 1.710 1.795 ;
        RECT  1.120 0.470 1.340 0.885 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.430 1.915 0.670 2.075 ;
    END
END AO31D1

MACRO AO31D2
    CLASS CORE ;
    FOREIGN AO31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.960 1.970 2.100 ;
        RECT  1.970 1.390 2.010 2.100 ;
        RECT  1.970 0.420 2.010 0.900 ;
        RECT  2.010 0.420 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.780 2.150 1.515 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.045 0.410 1.270 ;
        RECT  0.410 1.000 0.550 1.510 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.700 1.270 ;
        RECT  0.700 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.520 0.300 ;
        RECT  1.520 -0.300 1.740 0.340 ;
        RECT  1.740 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 1.915 1.450 2.075 ;
        RECT  0.670 1.915 1.210 2.050 ;
        RECT  1.710 0.765 1.850 1.795 ;
        RECT  1.340 0.765 1.710 0.885 ;
        RECT  0.260 1.635 1.710 1.795 ;
        RECT  1.120 0.470 1.340 0.885 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.430 1.915 0.670 2.075 ;
    END
END AO31D2

MACRO AO31D4
    CLASS CORE ;
    FOREIGN AO31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.780 1.650 4.110 2.030 ;
        RECT  3.780 0.490 4.110 0.870 ;
        RECT  4.110 0.490 4.530 2.030 ;
        RECT  4.530 1.650 4.690 2.030 ;
        RECT  4.530 0.490 4.690 0.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.710 1.330 1.340 ;
        RECT  1.330 0.710 2.970 0.830 ;
        RECT  2.970 0.710 3.120 1.235 ;
        RECT  3.120 0.950 3.170 1.110 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.480 0.950 1.690 1.110 ;
        RECT  1.690 0.950 1.830 1.515 ;
        RECT  1.830 1.395 2.590 1.515 ;
        RECT  2.590 1.130 2.750 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.000 0.560 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 0.980 0.300 ;
        RECT  0.980 -0.300 1.200 0.340 ;
        RECT  1.200 -0.300 2.900 0.300 ;
        RECT  2.900 -0.300 3.120 0.340 ;
        RECT  3.120 -0.300 3.370 0.300 ;
        RECT  3.370 -0.300 3.590 0.340 ;
        RECT  3.590 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 1.930 3.370 2.090 ;
        RECT  2.590 1.930 3.130 2.050 ;
        RECT  2.370 1.930 2.590 2.090 ;
        RECT  1.830 1.930 2.370 2.050 ;
        RECT  1.610 1.930 1.830 2.090 ;
        RECT  1.070 1.930 1.610 2.050 ;
        RECT  0.850 1.630 1.070 2.050 ;
        RECT  0.290 1.930 0.850 2.050 ;
        RECT  3.610 1.080 3.890 1.240 ;
        RECT  3.490 0.470 3.610 1.810 ;
        RECT  2.210 0.470 3.490 0.590 ;
        RECT  1.210 1.650 3.490 1.810 ;
        RECT  1.990 0.430 2.210 0.590 ;
        RECT  0.780 0.470 1.990 0.590 ;
        RECT  0.560 0.430 0.780 0.850 ;
        RECT  0.070 1.630 0.290 2.050 ;
        LAYER M1 ;
        RECT  3.780 0.490 3.895 0.870 ;
        RECT  3.780 1.650 3.895 2.030 ;
    END
END AO31D4

MACRO AO32D0
    CLASS CORE ;
    FOREIGN AO32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.660 2.790 1.710 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.985 1.830 1.515 ;
        RECT  1.830 0.985 1.870 1.225 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.985 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.230 1.515 ;
        RECT  0.230 0.985 0.260 1.225 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.985 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 1.840 0.300 ;
        RECT  1.840 -0.300 2.060 0.340 ;
        RECT  2.060 -0.300 2.250 0.300 ;
        RECT  2.250 -0.300 2.470 0.340 ;
        RECT  2.470 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.310 2.820 ;
        RECT  2.310 2.180 2.530 2.820 ;
        RECT  2.530 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 1.880 2.190 2.050 ;
        RECT  1.430 1.930 1.950 2.050 ;
        RECT  1.210 1.880 1.430 2.050 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.300 0.470 2.460 1.760 ;
        RECT  1.130 0.470 2.300 0.630 ;
        RECT  1.050 1.640 2.300 1.760 ;
        RECT  0.830 1.640 1.050 1.810 ;
        RECT  0.260 1.640 0.830 1.760 ;
        RECT  0.430 1.880 0.670 2.050 ;
        RECT  0.100 1.640 0.260 1.980 ;
    END
END AO32D0

MACRO AO32D1
    CLASS CORE ;
    FOREIGN AO32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.910 1.930 2.150 2.090 ;
        RECT  1.430 1.930 1.910 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.350 0.765 2.510 1.810 ;
        RECT  1.370 0.765 2.350 0.885 ;
        RECT  0.260 1.650 2.350 1.810 ;
        RECT  1.150 0.470 1.370 0.885 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AO32D1

MACRO AO32D2
    CLASS CORE ;
    FOREIGN AO32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.960 2.590 2.100 ;
        RECT  2.590 1.390 2.650 2.100 ;
        RECT  2.590 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.750 2.100 ;
        RECT  2.750 1.960 2.780 2.100 ;
        RECT  2.750 0.780 2.790 1.515 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.910 1.930 2.150 2.090 ;
        RECT  1.430 1.930 1.910 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.310 0.765 2.470 1.810 ;
        RECT  1.370 0.765 2.310 0.885 ;
        RECT  0.260 1.650 2.310 1.810 ;
        RECT  1.150 0.470 1.370 0.885 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AO32D2

MACRO AO32D4
    CLASS CORE ;
    FOREIGN AO32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.390 1.650 4.750 2.030 ;
        RECT  4.390 0.490 4.750 0.870 ;
        RECT  4.750 0.490 5.170 2.030 ;
        RECT  5.170 1.650 5.320 2.030 ;
        RECT  5.170 0.490 5.320 0.870 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.260 1.515 ;
        RECT  1.260 1.030 1.420 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.710 1.850 1.255 ;
        RECT  1.850 0.710 3.460 0.830 ;
        RECT  3.460 0.710 3.620 1.190 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.950 2.150 1.515 ;
        RECT  2.150 0.950 2.200 1.170 ;
        RECT  2.150 1.395 3.120 1.515 ;
        RECT  3.120 1.150 3.280 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.440 0.300 ;
        RECT  1.440 -0.300 1.660 0.340 ;
        RECT  1.660 -0.300 3.590 0.300 ;
        RECT  3.590 -0.300 3.810 0.340 ;
        RECT  3.810 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.720 1.915 3.960 2.075 ;
        RECT  3.180 1.915 3.720 2.050 ;
        RECT  2.960 1.915 3.180 2.075 ;
        RECT  2.420 1.915 2.960 2.050 ;
        RECT  2.200 1.915 2.420 2.075 ;
        RECT  1.660 1.915 2.200 2.050 ;
        RECT  1.440 1.635 1.660 2.050 ;
        RECT  0.970 1.890 1.440 2.050 ;
        RECT  0.750 1.635 0.970 2.050 ;
        RECT  0.280 1.910 0.750 2.050 ;
        RECT  4.110 0.470 4.270 1.795 ;
        RECT  2.800 0.470 4.110 0.590 ;
        RECT  1.800 1.635 4.110 1.795 ;
        RECT  2.580 0.430 2.800 0.590 ;
        RECT  0.980 0.470 2.580 0.590 ;
        RECT  0.760 0.450 0.980 0.870 ;
        RECT  0.060 1.635 0.280 2.050 ;
        LAYER M1 ;
        RECT  4.390 0.490 4.535 0.870 ;
        RECT  4.390 1.650 4.535 2.030 ;
    END
END AO32D4

MACRO AO33D0
    CLASS CORE ;
    FOREIGN AO33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.440 2.790 1.790 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.725 2.170 1.255 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.255 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.530 1.255 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.255 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.345 ;
        RECT  2.390 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 1.680 1.730 2.820 ;
        RECT  1.730 2.220 2.240 2.820 ;
        RECT  2.240 2.180 2.460 2.820 ;
        RECT  2.460 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.485 2.510 1.560 ;
        RECT  1.360 0.485 2.350 0.605 ;
        RECT  1.010 1.440 2.350 1.560 ;
        RECT  1.120 0.445 1.360 0.605 ;
        RECT  0.070 1.580 0.890 1.740 ;
        RECT  0.890 1.440 1.010 1.740 ;
    END
END AO33D0

MACRO AO33D1
    CLASS CORE ;
    FOREIGN AO33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 1.390 2.660 2.100 ;
        RECT  2.630 0.420 2.660 0.955 ;
        RECT  2.660 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.260 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 1.930 2.140 2.090 ;
        RECT  1.430 1.930 1.900 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.460 1.050 2.540 1.270 ;
        RECT  2.340 0.765 2.460 1.810 ;
        RECT  1.350 0.765 2.340 0.885 ;
        RECT  0.290 1.650 2.340 1.810 ;
        RECT  1.130 0.470 1.350 0.885 ;
        RECT  0.070 1.650 0.290 2.070 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AO33D1

MACRO AO33D2
    CLASS CORE ;
    FOREIGN AO33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.960 2.730 2.100 ;
        RECT  2.630 0.420 2.790 0.905 ;
        RECT  2.730 1.390 2.890 2.100 ;
        RECT  2.890 1.960 2.920 2.100 ;
        RECT  2.890 1.390 2.970 1.515 ;
        RECT  2.790 0.785 2.970 0.905 ;
        RECT  2.970 0.785 3.110 1.515 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.260 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 3.015 0.300 ;
        RECT  3.015 -0.300 3.235 0.340 ;
        RECT  3.235 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.300 2.820 ;
        RECT  2.300 2.180 2.520 2.820 ;
        RECT  2.520 2.220 3.115 2.820 ;
        RECT  3.115 2.180 3.335 2.820 ;
        RECT  3.335 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 1.930 2.140 2.090 ;
        RECT  1.430 1.930 1.900 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.460 1.080 2.690 1.245 ;
        RECT  2.340 0.765 2.460 1.810 ;
        RECT  1.350 0.765 2.340 0.885 ;
        RECT  0.290 1.650 2.340 1.810 ;
        RECT  1.130 0.470 1.350 0.885 ;
        RECT  0.430 1.930 0.670 2.090 ;
        RECT  0.070 1.650 0.290 2.070 ;
    END
END AO33D2

MACRO AO33D4
    CLASS CORE ;
    FOREIGN AO33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.070 1.650 5.390 2.030 ;
        RECT  5.070 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.980 2.030 ;
        RECT  5.810 0.490 5.980 0.870 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 0.750 0.500 1.190 ;
        RECT  2.010 1.070 2.040 1.515 ;
        RECT  0.500 0.750 2.040 0.870 ;
        RECT  2.040 0.750 2.170 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.150 0.840 1.515 ;
        RECT  0.840 1.395 1.690 1.515 ;
        RECT  1.630 0.990 1.690 1.140 ;
        RECT  1.690 0.990 1.830 1.515 ;
        RECT  1.830 0.990 1.850 1.140 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.750 2.710 1.310 ;
        RECT  2.710 0.750 4.250 0.870 ;
        RECT  4.250 0.750 4.410 1.235 ;
        RECT  4.410 1.005 4.710 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.990 2.970 1.140 ;
        RECT  2.970 0.990 3.110 1.475 ;
        RECT  3.110 1.355 3.870 1.475 ;
        RECT  3.870 1.005 4.030 1.475 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 2.280 0.300 ;
        RECT  2.280 -0.300 2.500 0.340 ;
        RECT  2.500 -0.300 4.330 0.300 ;
        RECT  4.330 -0.300 4.550 0.340 ;
        RECT  4.550 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.370 1.890 4.670 2.050 ;
        RECT  2.150 1.635 2.370 2.050 ;
        RECT  1.680 1.890 2.150 2.050 ;
        RECT  1.460 1.635 1.680 2.050 ;
        RECT  0.970 1.890 1.460 2.050 ;
        RECT  0.750 1.635 0.970 2.050 ;
        RECT  0.280 1.890 0.750 2.050 ;
        RECT  4.950 1.080 5.175 1.240 ;
        RECT  4.830 0.470 4.950 1.770 ;
        RECT  1.110 0.470 4.830 0.630 ;
        RECT  2.510 1.610 4.830 1.770 ;
        RECT  0.060 1.630 0.280 2.050 ;
        LAYER M1 ;
        RECT  5.070 0.490 5.175 0.870 ;
        RECT  5.070 1.650 5.175 2.030 ;
    END
END AO33D4

MACRO AOI211D0
    CLASS CORE ;
    FOREIGN AOI211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.450 0.590 0.605 ;
        RECT  0.590 0.470 1.310 0.605 ;
        RECT  0.990 1.660 1.370 1.820 ;
        RECT  1.310 0.450 1.370 0.605 ;
        RECT  1.370 0.450 1.530 1.820 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.235 ;
        RECT  0.550 0.860 0.740 1.020 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.170 0.870 1.795 ;
        RECT  0.870 1.170 0.930 1.390 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.080 1.250 1.300 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.600 2.820 ;
        END
    END VDD
END AOI211D0

MACRO AOI211D1
    CLASS CORE ;
    FOREIGN AOI211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 0.450 0.730 0.870 ;
        RECT  0.730 0.750 1.540 0.870 ;
        RECT  1.230 1.640 1.690 1.800 ;
        RECT  1.540 0.450 1.690 0.870 ;
        RECT  1.690 0.450 1.760 1.800 ;
        RECT  1.760 0.750 1.830 1.800 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.570 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 0.900 0.300 ;
        RECT  0.900 -0.300 1.120 0.340 ;
        RECT  1.120 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.200 2.820 ;
        RECT  0.200 2.180 0.420 2.820 ;
        RECT  0.420 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.630 1.920 1.850 2.080 ;
        RECT  1.090 1.920 1.630 2.040 ;
        RECT  0.870 1.660 1.090 2.080 ;
    END
END AOI211D1

MACRO AOI211D2
    CLASS CORE ;
    FOREIGN AOI211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.430 0.650 0.590 ;
        RECT  0.650 0.470 1.140 0.590 ;
        RECT  1.140 0.430 1.360 0.590 ;
        RECT  1.360 0.470 2.150 0.590 ;
        RECT  2.150 0.430 2.370 0.590 ;
        RECT  1.750 1.590 2.970 1.750 ;
        RECT  2.370 0.470 2.970 0.590 ;
        RECT  2.970 0.470 3.110 1.750 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.270 ;
        RECT  0.250 0.725 1.280 0.845 ;
        RECT  1.280 0.725 1.440 1.270 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.725 1.840 1.290 ;
        RECT  1.840 0.725 2.690 0.845 ;
        RECT  2.690 0.725 2.850 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.810 0.300 ;
        RECT  2.810 -0.300 3.030 0.340 ;
        RECT  3.030 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.730 2.820 ;
        RECT  0.730 2.180 0.950 2.820 ;
        RECT  0.950 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.420 1.390 1.580 2.100 ;
        RECT  1.580 1.890 1.610 2.100 ;
        RECT  1.610 1.890 3.130 2.050 ;
        RECT  1.390 1.915 1.420 2.100 ;
        RECT  0.290 1.915 1.390 2.050 ;
        RECT  0.260 1.915 0.290 2.100 ;
        RECT  0.100 1.390 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
    END
END AOI211D2

MACRO AOI211D4
    CLASS CORE ;
    FOREIGN AOI211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  1.625 1.430 1.845 1.810 ;
        RECT  1.845 1.430 1.870 1.550 ;
        RECT  0.430 0.710 1.870 0.870 ;
        RECT  1.870 0.710 2.290 1.550 ;
        RECT  2.290 1.430 2.385 1.550 ;
        RECT  2.385 1.430 2.605 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  2.290 0.710 3.790 0.870 ;
        RECT  3.790 0.450 4.010 0.870 ;
        RECT  4.010 0.750 4.480 0.870 ;
        RECT  4.480 0.450 4.700 0.870 ;
        RECT  4.700 0.750 5.280 0.870 ;
        RECT  5.280 0.450 5.500 0.870 ;
        RECT  5.500 0.750 5.970 0.870 ;
        RECT  5.970 0.450 6.190 0.870 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.390 0.300 ;
        RECT  3.390 -0.300 3.610 0.340 ;
        RECT  3.610 -0.300 4.880 0.300 ;
        RECT  4.880 -0.300 5.100 0.340 ;
        RECT  5.100 -0.300 6.370 0.300 ;
        RECT  6.370 -0.300 6.590 0.340 ;
        RECT  6.590 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.470 3.230 0.590 ;
        RECT  4.630 1.670 4.850 2.050 ;
        RECT  4.090 1.930 4.630 2.050 ;
        RECT  3.870 1.670 4.090 2.050 ;
        RECT  2.985 1.930 3.870 2.050 ;
        RECT  2.765 1.670 2.985 2.050 ;
        RECT  2.225 1.930 2.765 2.050 ;
        RECT  2.005 1.670 2.225 2.050 ;
        RECT  1.465 1.930 2.005 2.050 ;
        RECT  1.245 1.670 1.465 2.050 ;
        RECT  0.705 1.930 1.245 2.050 ;
        RECT  6.390 1.430 6.610 1.830 ;
        RECT  5.920 1.430 6.390 1.550 ;
        RECT  5.700 1.430 5.920 1.830 ;
        RECT  5.230 1.430 5.700 1.550 ;
        RECT  5.010 1.430 5.230 1.830 ;
        RECT  4.470 1.430 5.010 1.550 ;
        RECT  4.250 1.430 4.470 1.810 ;
        RECT  3.710 1.430 4.250 1.550 ;
        RECT  3.490 1.430 3.710 1.810 ;
        RECT  0.485 1.670 0.705 2.050 ;
        RECT  0.070 0.470 0.290 0.890 ;
        LAYER M1 ;
        RECT  0.430 0.710 1.655 0.870 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  1.625 1.430 1.655 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  3.790 0.450 4.010 0.870 ;
        RECT  4.010 0.750 4.480 0.870 ;
        RECT  4.480 0.450 4.700 0.870 ;
        RECT  4.700 0.750 5.280 0.870 ;
        RECT  5.280 0.450 5.500 0.870 ;
        RECT  5.500 0.750 5.970 0.870 ;
        RECT  5.970 0.450 6.190 0.870 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  2.505 1.430 2.605 1.810 ;
        RECT  2.505 0.710 3.790 0.870 ;
    END
END AOI211D4

MACRO AOI21D0
    CLASS CORE ;
    FOREIGN AOI21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.470 0.560 1.740 ;
        RECT  0.560 0.470 0.660 0.600 ;
        RECT  0.660 0.440 0.900 0.600 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 0.920 0.710 1.140 ;
        RECT  0.710 0.725 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.280 2.820 ;
        END
    END VDD
END AOI21D0

MACRO AOI21D1
    CLASS CORE ;
    FOREIGN AOI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.795 ;
        RECT  0.550 1.635 0.730 1.795 ;
        RECT  0.550 0.725 0.790 0.870 ;
        RECT  0.790 0.450 1.010 0.870 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.200 0.300 ;
        RECT  1.200 -0.300 1.420 0.340 ;
        RECT  1.420 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.260 2.820 ;
        RECT  1.260 2.180 1.480 2.820 ;
        RECT  1.480 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.870 1.635 1.090 2.050 ;
        RECT  0.330 1.930 0.870 2.050 ;
        RECT  0.090 1.930 0.330 2.090 ;
    END
END AOI21D1

MACRO AOI21D2
    CLASS CORE ;
    FOREIGN AOI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 0.470 0.500 0.605 ;
        RECT  0.500 0.470 0.660 1.125 ;
        RECT  0.660 1.005 0.730 1.125 ;
        RECT  0.730 1.005 0.870 1.770 ;
        RECT  0.660 0.470 1.520 0.605 ;
        RECT  1.520 0.445 1.760 0.605 ;
        RECT  0.870 1.610 2.130 1.770 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.260 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.725 1.200 1.290 ;
        RECT  1.200 0.725 2.010 0.845 ;
        RECT  2.010 0.725 2.150 1.290 ;
        RECT  2.150 1.050 2.190 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.870 0.300 ;
        RECT  0.870 -0.300 1.090 0.340 ;
        RECT  1.090 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.460 1.960 2.490 2.100 ;
        RECT  2.300 1.370 2.460 2.100 ;
        RECT  2.270 1.890 2.300 2.100 ;
        RECT  0.280 1.890 2.270 2.050 ;
        RECT  0.060 1.640 0.280 2.070 ;
    END
END AOI21D2

MACRO AOI21D4
    CLASS CORE ;
    FOREIGN AOI21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  1.625 1.430 1.845 1.810 ;
        RECT  1.845 1.430 1.870 1.550 ;
        RECT  0.430 0.710 1.870 0.870 ;
        RECT  1.870 0.710 2.290 1.550 ;
        RECT  2.290 1.430 2.385 1.550 ;
        RECT  2.385 1.430 2.605 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  2.290 0.710 3.790 0.850 ;
        RECT  3.790 0.430 4.010 0.850 ;
        RECT  4.010 0.710 4.480 0.850 ;
        RECT  4.480 0.430 4.700 0.850 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.390 0.300 ;
        RECT  3.390 -0.300 3.610 0.340 ;
        RECT  3.610 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.470 3.230 0.590 ;
        RECT  4.480 1.630 4.700 2.050 ;
        RECT  4.010 1.890 4.480 2.050 ;
        RECT  3.790 1.630 4.010 2.050 ;
        RECT  2.985 1.930 3.790 2.050 ;
        RECT  2.765 1.670 2.985 2.050 ;
        RECT  2.225 1.930 2.765 2.050 ;
        RECT  2.005 1.670 2.225 2.050 ;
        RECT  1.465 1.930 2.005 2.050 ;
        RECT  1.245 1.670 1.465 2.050 ;
        RECT  0.705 1.930 1.245 2.050 ;
        RECT  0.070 0.470 0.290 0.890 ;
        RECT  0.485 1.670 0.705 2.050 ;
        LAYER M1 ;
        RECT  3.790 0.430 4.010 0.850 ;
        RECT  4.010 0.710 4.480 0.850 ;
        RECT  4.480 0.430 4.700 0.850 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  1.625 1.430 1.655 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.430 0.710 1.655 0.870 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  2.505 1.430 2.605 1.810 ;
        RECT  2.505 0.710 3.790 0.850 ;
    END
END AOI21D4

MACRO AOI221D0
    CLASS CORE ;
    FOREIGN AOI221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.440 0.550 1.495 ;
        RECT  0.550 0.440 0.700 0.600 ;
        RECT  0.550 1.375 0.900 1.495 ;
        RECT  0.900 1.375 1.020 1.810 ;
        RECT  1.020 1.650 1.440 1.810 ;
        RECT  0.700 0.470 1.810 0.600 ;
        RECT  1.810 0.440 2.050 0.600 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END C
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.725 0.870 1.255 ;
        RECT  0.870 1.015 0.880 1.255 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.980 1.830 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 0.720 1.210 0.880 ;
        RECT  1.210 0.720 2.000 0.860 ;
        RECT  2.000 0.720 2.160 1.255 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.660 1.930 1.980 2.050 ;
        RECT  1.980 1.600 2.140 2.050 ;
        RECT  0.500 1.620 0.660 2.050 ;
    END
END AOI221D0

MACRO AOI221D1
    CLASS CORE ;
    FOREIGN AOI221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 0.465 0.690 0.885 ;
        RECT  0.690 0.765 1.510 0.885 ;
        RECT  1.510 0.465 1.730 0.885 ;
        RECT  1.880 1.650 2.330 1.810 ;
        RECT  1.730 0.765 2.330 0.885 ;
        RECT  2.330 0.765 2.470 1.810 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.130 0.300 ;
        RECT  1.130 -0.300 1.350 0.340 ;
        RECT  1.350 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.340 ;
        RECT  2.390 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.180 1.930 1.400 2.090 ;
        RECT  0.640 1.930 1.180 2.050 ;
        RECT  0.610 1.930 0.640 2.090 ;
        RECT  0.450 1.360 0.610 2.090 ;
        RECT  2.280 1.930 2.500 2.090 ;
        RECT  1.740 1.930 2.280 2.050 ;
        RECT  1.520 1.650 1.740 2.070 ;
        RECT  0.780 1.650 1.520 1.810 ;
        RECT  0.420 1.950 0.450 2.090 ;
    END
END AOI221D1

MACRO AOI221D2
    CLASS CORE ;
    FOREIGN AOI221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.470 0.290 0.885 ;
        RECT  0.290 0.765 0.870 0.885 ;
        RECT  0.870 0.470 1.090 0.885 ;
        RECT  1.090 0.765 2.200 0.885 ;
        RECT  2.200 0.470 2.425 0.885 ;
        RECT  2.425 0.765 2.650 0.885 ;
        RECT  2.650 0.765 2.790 1.810 ;
        RECT  2.790 0.470 3.015 0.885 ;
        RECT  3.015 0.765 4.120 0.885 ;
        RECT  2.790 1.650 4.190 1.810 ;
        RECT  4.120 0.470 4.340 0.885 ;
        RECT  4.190 1.650 4.410 2.070 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.070 1.235 ;
        RECT  1.070 1.005 1.190 1.515 ;
        RECT  1.190 1.395 2.080 1.515 ;
        RECT  2.080 1.030 2.240 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.005 3.110 1.515 ;
        RECT  3.110 1.395 4.000 1.515 ;
        RECT  4.000 1.030 4.160 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.540 0.300 ;
        RECT  1.540 -0.300 1.760 0.340 ;
        RECT  1.760 -0.300 3.450 0.300 ;
        RECT  3.450 -0.300 3.670 0.340 ;
        RECT  3.670 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 1.930 1.930 2.050 ;
        RECT  1.930 1.930 2.150 2.090 ;
        RECT  2.150 1.930 3.050 2.050 ;
        RECT  3.050 1.930 3.270 2.090 ;
        RECT  3.270 1.930 3.810 2.050 ;
        RECT  3.810 1.930 4.050 2.090 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.260 1.650 0.790 1.790 ;
        RECT  0.790 1.650 1.010 2.070 ;
        RECT  1.010 1.650 2.530 1.810 ;
        RECT  1.150 1.930 1.390 2.090 ;
        RECT  0.070 1.960 0.100 2.100 ;
    END
END AOI221D2

MACRO AOI221D4
    CLASS CORE ;
    FOREIGN AOI221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.640 2.830 2.020 ;
        RECT  2.590 0.760 2.830 0.920 ;
        RECT  2.830 0.760 3.250 2.020 ;
        RECT  3.250 0.760 3.620 0.920 ;
        RECT  3.250 1.640 3.670 2.020 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.160 0.300 ;
        RECT  1.160 -0.300 1.380 0.340 ;
        RECT  1.380 -0.300 2.220 0.300 ;
        RECT  2.220 -0.300 2.440 0.340 ;
        RECT  2.440 -0.300 3.000 0.300 ;
        RECT  3.000 -0.300 3.220 0.340 ;
        RECT  3.220 -0.300 3.790 0.300 ;
        RECT  3.790 -0.300 4.010 0.340 ;
        RECT  4.010 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 1.930 1.980 2.100 ;
        RECT  1.980 1.370 2.140 2.100 ;
        RECT  2.140 1.960 2.170 2.100 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  0.830 1.640 1.050 2.050 ;
        RECT  1.050 1.640 1.810 1.800 ;
        RECT  1.410 1.930 1.950 2.050 ;
        RECT  4.100 1.050 4.140 1.270 ;
        RECT  3.980 0.470 4.100 1.270 ;
        RECT  2.040 0.470 3.980 0.590 ;
        RECT  1.820 0.470 2.040 0.885 ;
        RECT  1.000 0.765 1.820 0.885 ;
        RECT  0.780 0.470 1.000 0.885 ;
        RECT  0.540 0.765 0.780 0.885 ;
        RECT  0.540 1.640 0.690 1.800 ;
        RECT  4.380 1.960 4.410 2.100 ;
        RECT  4.260 0.420 4.380 2.100 ;
        RECT  4.220 0.420 4.260 0.900 ;
        RECT  4.220 1.390 4.260 2.100 ;
        RECT  3.760 1.390 4.220 1.510 ;
        RECT  4.190 1.960 4.220 2.100 ;
        RECT  0.420 0.765 0.540 1.800 ;
        RECT  1.170 1.930 1.410 2.090 ;
        RECT  0.070 1.635 0.290 2.050 ;
        RECT  3.600 1.050 3.760 1.510 ;
        LAYER M1 ;
        RECT  3.465 1.640 3.670 2.020 ;
        RECT  3.465 0.760 3.620 0.920 ;
        RECT  2.590 0.760 2.615 0.920 ;
    END
END AOI221D4

MACRO AOI222D0
    CLASS CORE ;
    FOREIGN AOI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.430 0.870 1.510 ;
        RECT  0.870 0.430 1.020 0.590 ;
        RECT  0.870 1.390 1.520 1.510 ;
        RECT  1.520 1.390 1.640 1.810 ;
        RECT  1.640 1.650 1.760 1.810 ;
        RECT  1.020 0.470 2.120 0.590 ;
        RECT  2.120 0.430 2.360 0.590 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.570 1.235 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 0.720 1.530 0.880 ;
        RECT  1.530 0.720 2.310 0.840 ;
        RECT  2.310 0.720 2.470 1.255 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.270 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.960 2.150 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.460 0.300 ;
        RECT  1.460 -0.300 1.680 0.340 ;
        RECT  1.680 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.430 2.820 ;
        RECT  0.430 2.180 0.650 2.820 ;
        RECT  0.650 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.980 1.930 2.300 2.050 ;
        RECT  2.300 1.600 2.460 2.050 ;
        RECT  0.820 1.630 0.980 2.050 ;
        RECT  0.260 1.930 0.820 2.050 ;
        RECT  0.100 1.610 0.260 2.050 ;
    END
END AOI222D0

MACRO AOI222D1
    CLASS CORE ;
    FOREIGN AOI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 0.470 1.010 0.885 ;
        RECT  1.010 0.765 1.850 0.885 ;
        RECT  1.850 0.470 2.070 0.885 ;
        RECT  2.190 1.410 2.330 1.810 ;
        RECT  2.070 0.765 2.330 0.885 ;
        RECT  2.330 0.765 2.410 1.810 ;
        RECT  2.410 0.765 2.470 1.550 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.490 0.300 ;
        RECT  1.490 -0.300 1.710 0.340 ;
        RECT  1.710 -0.300 2.510 0.300 ;
        RECT  2.510 -0.300 2.730 0.340 ;
        RECT  2.730 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 1.930 1.540 2.050 ;
        RECT  1.540 1.930 1.760 2.090 ;
        RECT  0.780 1.635 1.000 2.050 ;
        RECT  0.290 1.930 0.780 2.050 ;
        RECT  0.260 1.930 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  2.570 1.650 2.790 2.070 ;
        RECT  2.000 1.930 2.570 2.050 ;
        RECT  1.880 1.360 2.000 2.050 ;
        RECT  1.840 1.360 1.880 1.810 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  1.140 1.650 1.840 1.810 ;
    END
END AOI222D1

MACRO AOI222D2
    CLASS CORE ;
    FOREIGN AOI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 0.470 1.020 0.885 ;
        RECT  1.020 0.765 2.200 0.885 ;
        RECT  2.200 0.470 2.420 0.885 ;
        RECT  2.420 0.765 4.060 0.885 ;
        RECT  4.060 0.470 4.280 0.885 ;
        RECT  4.840 1.960 4.870 2.100 ;
        RECT  3.300 1.640 4.870 1.800 ;
        RECT  4.280 0.765 4.870 0.885 ;
        RECT  4.870 0.765 5.030 2.100 ;
        RECT  5.030 1.960 5.060 2.100 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.520 ;
        RECT  0.250 1.400 1.350 1.520 ;
        RECT  1.350 1.030 1.510 1.520 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.030 1.860 1.520 ;
        RECT  1.860 1.400 2.650 1.520 ;
        RECT  2.650 1.005 2.770 1.520 ;
        RECT  2.770 1.005 3.110 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.590 1.235 ;
        RECT  3.590 1.005 3.750 1.520 ;
        RECT  3.750 1.400 4.570 1.520 ;
        RECT  4.570 1.030 4.730 1.520 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.490 0.300 ;
        RECT  1.490 -0.300 1.710 0.340 ;
        RECT  1.710 -0.300 2.860 0.300 ;
        RECT  2.860 -0.300 3.080 0.340 ;
        RECT  3.080 -0.300 3.400 0.300 ;
        RECT  3.400 -0.300 3.620 0.340 ;
        RECT  3.620 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.940 0.340 ;
        RECT  4.940 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.660 1.640 3.180 1.800 ;
        RECT  1.440 1.640 1.660 2.070 ;
        RECT  0.970 1.640 1.440 1.780 ;
        RECT  0.750 1.640 0.970 2.070 ;
        RECT  0.280 1.640 0.750 1.780 ;
        RECT  4.440 1.930 4.680 2.090 ;
        RECT  3.900 1.930 4.440 2.050 ;
        RECT  3.680 1.930 3.900 2.090 ;
        RECT  2.800 1.930 3.680 2.050 ;
        RECT  2.580 1.930 2.800 2.090 ;
        RECT  2.040 1.930 2.580 2.050 ;
        RECT  0.060 1.640 0.280 2.070 ;
        RECT  1.800 1.930 2.040 2.090 ;
    END
END AOI222D2

MACRO AOI222D4
    CLASS CORE ;
    FOREIGN AOI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.030 1.640 3.150 2.020 ;
        RECT  2.930 0.760 3.150 0.920 ;
        RECT  3.150 0.760 3.570 2.020 ;
        RECT  3.570 0.760 3.950 0.920 ;
        RECT  3.570 1.640 3.990 2.020 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.725 1.210 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.530 1.270 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.830 0.300 ;
        RECT  0.830 -0.300 1.050 0.340 ;
        RECT  1.050 -0.300 2.560 0.300 ;
        RECT  2.560 -0.300 2.780 0.340 ;
        RECT  2.780 -0.300 3.340 0.300 ;
        RECT  3.340 -0.300 3.560 0.340 ;
        RECT  3.560 -0.300 4.120 0.300 ;
        RECT  4.120 -0.300 4.340 0.340 ;
        RECT  4.340 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.770 0.470 0.890 0.885 ;
        RECT  0.890 0.470 1.500 0.590 ;
        RECT  1.500 0.430 1.720 0.590 ;
        RECT  1.720 0.470 1.920 0.590 ;
        RECT  1.920 0.470 2.140 0.885 ;
        RECT  2.140 0.470 4.270 0.590 ;
        RECT  4.270 0.470 4.420 1.270 ;
        RECT  4.420 1.050 4.430 1.270 ;
        RECT  1.430 1.400 2.290 1.540 ;
        RECT  2.290 1.400 2.510 2.080 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  0.830 1.640 1.050 2.090 ;
        RECT  1.050 1.930 1.590 2.050 ;
        RECT  1.590 1.660 1.810 2.090 ;
        RECT  0.570 0.765 0.770 0.885 ;
        RECT  0.570 1.640 0.690 1.800 ;
        RECT  0.450 0.765 0.570 1.800 ;
        RECT  0.390 0.765 0.450 0.885 ;
        RECT  4.700 1.960 4.730 2.100 ;
        RECT  4.560 0.420 4.700 2.100 ;
        RECT  4.540 0.420 4.560 0.900 ;
        RECT  4.540 1.390 4.560 2.100 ;
        RECT  4.080 1.390 4.540 1.510 ;
        RECT  4.510 1.960 4.540 2.100 ;
        RECT  0.170 0.470 0.390 0.885 ;
        RECT  1.210 1.400 1.430 1.810 ;
        RECT  3.920 1.050 4.080 1.510 ;
        RECT  0.070 1.640 0.290 2.090 ;
        LAYER M1 ;
        RECT  3.785 1.640 3.990 2.020 ;
        RECT  3.785 0.760 3.950 0.920 ;
    END
END AOI222D4

MACRO AOI22D0
    CLASS CORE ;
    FOREIGN AOI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.285 0.750 1.815 ;
        RECT  0.750 0.710 0.870 1.815 ;
        RECT  0.870 0.710 0.990 0.850 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 0.470 0.630 1.010 ;
        RECT  0.630 0.470 1.350 0.590 ;
        RECT  1.350 0.470 1.510 1.730 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.130 0.570 1.795 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.600 2.820 ;
        END
    END VDD
END AOI22D0

MACRO AOI22D1
    CLASS CORE ;
    FOREIGN AOI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.430 0.390 0.845 ;
        RECT  0.390 0.725 1.510 0.845 ;
        RECT  1.240 1.650 1.690 1.810 ;
        RECT  1.510 0.430 1.690 0.845 ;
        RECT  1.690 0.430 1.730 1.810 ;
        RECT  1.730 0.725 1.830 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.540 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.840 0.300 ;
        RECT  0.840 -0.300 1.060 0.340 ;
        RECT  1.060 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.280 1.930 0.880 2.050 ;
        RECT  0.880 1.635 1.100 2.050 ;
        RECT  1.100 1.930 1.640 2.050 ;
        RECT  1.640 1.930 1.860 2.090 ;
        RECT  0.060 1.635 0.280 2.050 ;
    END
END AOI22D1

MACRO AOI22D2
    CLASS CORE ;
    FOREIGN AOI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.430 1.100 0.590 ;
        RECT  1.100 0.470 1.690 0.590 ;
        RECT  1.690 0.470 1.830 1.530 ;
        RECT  1.830 1.410 2.060 1.530 ;
        RECT  2.060 1.410 2.280 1.810 ;
        RECT  1.830 0.470 2.440 0.590 ;
        RECT  2.440 0.430 2.680 0.590 ;
        RECT  2.280 1.410 2.820 1.530 ;
        RECT  2.820 1.410 3.040 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.725 0.550 1.290 ;
        RECT  0.550 0.725 1.410 0.845 ;
        RECT  1.410 0.725 1.570 1.290 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 0.725 2.160 1.290 ;
        RECT  2.160 0.725 2.970 0.845 ;
        RECT  2.970 0.725 3.130 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.220 0.300 ;
        RECT  0.220 -0.300 0.440 0.340 ;
        RECT  0.440 -0.300 1.670 0.300 ;
        RECT  1.670 -0.300 1.890 0.340 ;
        RECT  1.890 -0.300 3.100 0.300 ;
        RECT  3.100 -0.300 3.320 0.340 ;
        RECT  3.320 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 1.280 2.820 ;
        RECT  1.280 2.180 1.500 2.820 ;
        RECT  1.500 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.910 1.370 1.070 2.100 ;
        RECT  1.070 1.930 1.100 2.100 ;
        RECT  1.100 1.930 1.680 2.050 ;
        RECT  1.680 1.650 1.900 2.070 ;
        RECT  1.900 1.930 2.440 2.050 ;
        RECT  2.440 1.650 2.660 2.070 ;
        RECT  2.660 1.930 3.200 2.050 ;
        RECT  3.200 1.930 3.230 2.100 ;
        RECT  3.230 1.370 3.390 2.100 ;
        RECT  3.390 1.960 3.420 2.100 ;
        RECT  0.880 1.930 0.910 2.100 ;
        RECT  0.300 1.930 0.880 2.050 ;
        RECT  0.270 1.930 0.300 2.100 ;
        RECT  0.110 1.370 0.270 2.100 ;
        RECT  0.080 1.960 0.110 2.100 ;
    END
END AOI22D2

MACRO AOI22D4
    CLASS CORE ;
    FOREIGN AOI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  1.625 1.430 1.845 1.810 ;
        RECT  1.845 1.430 1.870 1.550 ;
        RECT  0.430 0.710 1.870 0.870 ;
        RECT  1.870 0.710 2.290 1.550 ;
        RECT  2.290 1.430 2.385 1.550 ;
        RECT  2.385 1.430 2.605 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  2.290 0.710 6.580 0.870 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.400 0.300 ;
        RECT  3.400 -0.300 3.620 0.340 ;
        RECT  3.620 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.505 2.820 ;
        RECT  3.505 2.180 3.725 2.820 ;
        RECT  3.725 2.220 4.300 2.820 ;
        RECT  4.300 2.180 4.520 2.820 ;
        RECT  4.520 2.220 5.090 2.820 ;
        RECT  5.090 2.180 5.310 2.820 ;
        RECT  5.310 2.220 5.890 2.820 ;
        RECT  5.890 2.180 6.110 2.820 ;
        RECT  6.110 2.220 6.690 2.820 ;
        RECT  6.690 2.180 6.910 2.820 ;
        RECT  6.910 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.470 3.240 0.590 ;
        RECT  6.290 1.630 6.510 2.050 ;
        RECT  5.710 1.890 6.290 2.050 ;
        RECT  5.490 1.630 5.710 2.050 ;
        RECT  4.910 1.890 5.490 2.050 ;
        RECT  4.690 1.630 4.910 2.050 ;
        RECT  4.125 1.890 4.690 2.050 ;
        RECT  3.905 1.630 4.125 2.050 ;
        RECT  2.985 1.930 3.905 2.050 ;
        RECT  2.765 1.670 2.985 2.050 ;
        RECT  2.225 1.930 2.765 2.050 ;
        RECT  2.005 1.670 2.225 2.050 ;
        RECT  1.465 1.930 2.005 2.050 ;
        RECT  1.245 1.670 1.465 2.050 ;
        RECT  0.705 1.930 1.245 2.050 ;
        RECT  6.720 0.470 6.940 0.890 ;
        RECT  0.485 1.670 0.705 2.050 ;
        RECT  0.070 0.470 0.290 0.890 ;
        RECT  3.780 0.470 6.720 0.590 ;
        LAYER M1 ;
        RECT  3.145 1.430 3.365 1.810 ;
        RECT  2.605 1.430 3.145 1.550 ;
        RECT  1.625 1.430 1.655 1.810 ;
        RECT  1.085 1.430 1.625 1.550 ;
        RECT  0.865 1.430 1.085 1.810 ;
        RECT  0.325 1.430 0.865 1.550 ;
        RECT  0.430 0.710 1.655 0.870 ;
        RECT  0.105 1.430 0.325 1.830 ;
        RECT  2.505 0.710 6.580 0.870 ;
        RECT  2.505 1.430 2.605 1.810 ;
    END
END AOI22D4

MACRO AOI31D0
    CLASS CORE ;
    FOREIGN AOI31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 1.640 0.260 1.980 ;
        RECT  0.260 1.640 0.830 1.760 ;
        RECT  0.830 1.640 1.050 1.810 ;
        RECT  1.050 1.640 1.690 1.760 ;
        RECT  1.110 0.470 1.690 0.630 ;
        RECT  1.690 0.470 1.830 1.760 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.540 0.300 ;
        RECT  1.540 -0.300 1.760 0.340 ;
        RECT  1.760 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 1.880 1.450 2.050 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.880 0.670 2.050 ;
    END
END AOI31D0

MACRO AOI31D1
    CLASS CORE ;
    FOREIGN AOI31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  1.130 0.470 1.350 0.885 ;
        RECT  0.260 1.650 1.690 1.810 ;
        RECT  1.350 0.765 1.690 0.885 ;
        RECT  1.690 0.765 1.830 1.810 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.530 1.270 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.160 0.300 ;
        RECT  0.160 -0.300 0.380 0.340 ;
        RECT  0.380 -0.300 1.540 0.300 ;
        RECT  1.540 -0.300 1.760 0.340 ;
        RECT  1.760 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 1.930 1.450 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AOI31D1

MACRO AOI31D2
    CLASS CORE ;
    FOREIGN AOI31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 0.430 0.860 0.850 ;
        RECT  0.860 0.470 2.105 0.590 ;
        RECT  2.105 0.430 2.325 0.590 ;
        RECT  1.310 1.640 3.290 1.800 ;
        RECT  2.325 0.470 3.290 0.590 ;
        RECT  3.290 0.470 3.430 1.800 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.990 0.570 1.515 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.390 1.235 ;
        RECT  1.390 1.005 1.510 1.515 ;
        RECT  1.510 1.395 3.010 1.515 ;
        RECT  3.010 0.910 3.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 0.725 1.790 1.170 ;
        RECT  1.790 0.725 2.650 0.845 ;
        RECT  2.650 0.725 2.810 1.255 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.230 0.300 ;
        RECT  0.230 -0.300 0.450 0.340 ;
        RECT  0.450 -0.300 1.050 0.300 ;
        RECT  1.050 -0.300 1.270 0.340 ;
        RECT  1.270 -0.300 3.150 0.300 ;
        RECT  3.150 -0.300 3.370 0.340 ;
        RECT  3.370 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.530 2.820 ;
        RECT  0.530 2.180 0.750 2.820 ;
        RECT  0.750 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 1.930 3.450 2.090 ;
        RECT  2.690 1.930 3.230 2.050 ;
        RECT  2.470 1.930 2.690 2.090 ;
        RECT  1.930 1.930 2.470 2.050 ;
        RECT  1.710 1.930 1.930 2.090 ;
        RECT  1.170 1.930 1.710 2.050 ;
        RECT  0.950 1.630 1.170 2.050 ;
        RECT  0.340 1.920 0.950 2.050 ;
        RECT  0.120 1.630 0.340 2.050 ;
    END
END AOI31D2

MACRO AOI31D4
    CLASS CORE ;
    FOREIGN AOI31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.145 1.650 0.365 2.050 ;
        RECT  0.470 0.710 1.620 0.830 ;
        RECT  1.620 0.710 1.740 1.070 ;
        RECT  0.365 1.650 3.790 1.770 ;
        RECT  1.740 0.950 3.790 1.070 ;
        RECT  3.790 0.950 4.090 1.770 ;
        RECT  4.090 0.750 4.210 1.770 ;
        RECT  4.210 1.650 5.305 1.770 ;
        RECT  4.210 0.750 5.710 0.870 ;
        RECT  5.710 0.450 5.930 0.870 ;
        RECT  5.930 0.750 6.400 0.870 ;
        RECT  6.400 0.450 6.620 0.870 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.825 1.325 2.010 1.485 ;
        RECT  2.010 1.285 2.470 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.310 0.300 ;
        RECT  5.310 -0.300 5.530 0.340 ;
        RECT  5.530 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.330 0.470 3.370 0.590 ;
        RECT  3.900 0.470 5.150 0.590 ;
        RECT  3.780 0.470 3.900 0.830 ;
        RECT  6.400 1.630 6.620 2.050 ;
        RECT  5.930 1.890 6.400 2.050 ;
        RECT  5.710 1.630 5.930 2.050 ;
        RECT  0.505 1.890 5.710 2.050 ;
        RECT  1.970 0.710 3.780 0.830 ;
        RECT  0.110 0.470 0.330 0.890 ;
        LAYER M1 ;
        RECT  6.400 0.450 6.620 0.870 ;
        RECT  5.930 0.750 6.400 0.870 ;
        RECT  5.710 0.450 5.930 0.870 ;
        RECT  1.740 0.950 3.575 1.070 ;
        RECT  1.620 0.710 1.740 1.070 ;
        RECT  0.365 1.650 3.575 1.770 ;
        RECT  0.145 1.650 0.365 2.050 ;
        RECT  0.470 0.710 1.620 0.830 ;
        RECT  4.425 1.650 5.305 1.770 ;
        RECT  4.425 0.750 5.710 0.870 ;
    END
END AOI31D4

MACRO AOI32D0
    CLASS CORE ;
    FOREIGN AOI32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 1.670 0.260 2.005 ;
        RECT  0.260 1.670 2.010 1.810 ;
        RECT  1.180 0.470 2.010 0.630 ;
        RECT  2.010 0.470 2.150 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.005 1.890 1.225 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.990 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.985 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.985 1.190 1.515 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.985 1.530 1.515 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 1.860 0.300 ;
        RECT  1.860 -0.300 2.080 0.340 ;
        RECT  2.080 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 1.930 2.170 2.070 ;
        RECT  1.430 1.930 1.950 2.050 ;
        RECT  1.210 1.930 1.430 2.070 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.930 0.670 2.070 ;
    END
END AOI32D0

MACRO AOI32D1
    CLASS CORE ;
    FOREIGN AOI32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  1.150 0.470 1.370 0.885 ;
        RECT  0.260 1.650 2.010 1.810 ;
        RECT  1.370 0.765 2.010 0.885 ;
        RECT  2.010 0.765 2.150 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.890 1.270 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 1.860 0.300 ;
        RECT  1.860 -0.300 2.080 0.340 ;
        RECT  2.080 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.430 1.930 1.930 2.050 ;
        RECT  1.930 1.930 2.170 2.090 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AOI32D1

MACRO AOI32D2
    CLASS CORE ;
    FOREIGN AOI32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 0.430 1.050 0.850 ;
        RECT  1.050 0.470 2.745 0.590 ;
        RECT  2.745 0.430 2.965 0.590 ;
        RECT  1.950 1.600 3.930 1.760 ;
        RECT  2.965 0.470 3.930 0.590 ;
        RECT  3.930 0.470 4.070 1.760 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.990 0.550 1.515 ;
        RECT  0.550 1.380 1.340 1.515 ;
        RECT  1.340 0.990 1.500 1.515 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.475 ;
        RECT  2.150 1.355 3.610 1.475 ;
        RECT  3.610 0.930 3.750 1.475 ;
        RECT  3.750 0.930 3.800 1.150 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 0.930 2.330 1.150 ;
        RECT  2.330 0.725 2.470 1.235 ;
        RECT  2.470 0.725 3.290 0.845 ;
        RECT  3.290 0.725 3.450 1.170 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.170 0.300 ;
        RECT  0.170 -0.300 0.390 0.340 ;
        RECT  0.390 -0.300 1.620 0.300 ;
        RECT  1.620 -0.300 1.840 0.340 ;
        RECT  1.840 -0.300 3.800 0.300 ;
        RECT  3.800 -0.300 4.020 0.340 ;
        RECT  4.020 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.590 1.620 1.810 2.040 ;
        RECT  1.810 1.920 2.350 2.040 ;
        RECT  2.350 1.880 4.090 2.040 ;
        RECT  1.050 1.920 1.590 2.040 ;
        RECT  0.830 1.635 1.050 2.040 ;
        RECT  0.290 1.920 0.830 2.040 ;
        RECT  0.070 1.620 0.290 2.040 ;
    END
END AOI32D2

MACRO AOI32D4
    CLASS CORE ;
    FOREIGN AOI32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.640 3.470 2.020 ;
        RECT  2.970 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 3.970 2.020 ;
        RECT  3.890 0.500 3.970 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.850 0.300 ;
        RECT  1.850 -0.300 2.070 0.340 ;
        RECT  2.070 -0.300 2.580 0.300 ;
        RECT  2.580 -0.300 2.800 0.340 ;
        RECT  2.800 -0.300 3.360 0.300 ;
        RECT  3.360 -0.300 3.580 0.340 ;
        RECT  3.580 -0.300 4.140 0.300 ;
        RECT  4.140 -0.300 4.360 0.340 ;
        RECT  4.360 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.360 2.820 ;
        RECT  3.360 2.180 3.580 2.820 ;
        RECT  3.580 2.220 4.140 2.820 ;
        RECT  4.140 2.180 4.360 2.820 ;
        RECT  4.360 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 1.930 2.140 2.090 ;
        RECT  1.430 1.930 1.900 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  2.090 1.080 2.270 1.240 ;
        RECT  1.970 0.755 2.090 1.810 ;
        RECT  1.365 0.755 1.970 0.885 ;
        RECT  0.290 1.650 1.970 1.810 ;
        RECT  1.145 0.470 1.365 0.885 ;
        RECT  2.520 1.080 3.080 1.240 ;
        RECT  2.400 0.790 2.520 1.480 ;
        RECT  2.380 0.790 2.400 0.910 ;
        RECT  2.380 1.360 2.400 1.480 ;
        RECT  2.220 0.420 2.380 0.910 ;
        RECT  2.220 1.360 2.380 1.680 ;
        RECT  0.070 1.650 0.290 2.070 ;
        RECT  0.430 1.930 0.670 2.090 ;
        LAYER M1 ;
        RECT  2.970 0.500 3.255 0.880 ;
        RECT  2.970 1.640 3.255 2.020 ;
    END
END AOI32D4

MACRO AOI33D0
    CLASS CORE ;
    FOREIGN AOI33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 1.650 0.260 1.980 ;
        RECT  0.260 1.650 0.830 1.770 ;
        RECT  0.830 1.650 1.050 1.810 ;
        RECT  1.050 1.650 2.330 1.770 ;
        RECT  1.150 0.490 2.330 0.650 ;
        RECT  2.330 0.490 2.470 1.770 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.005 2.200 1.225 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.985 1.850 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.520 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.985 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.985 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.985 1.210 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 1.890 2.160 2.050 ;
        RECT  1.430 1.930 1.920 2.050 ;
        RECT  1.210 1.890 1.430 2.050 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.890 0.670 2.050 ;
    END
END AOI33D0

MACRO AOI33D1
    CLASS CORE ;
    FOREIGN AOI33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  1.130 0.470 1.350 0.885 ;
        RECT  0.260 1.650 2.330 1.810 ;
        RECT  1.350 0.765 2.330 0.885 ;
        RECT  2.330 0.765 2.470 1.810 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 1.930 2.160 2.090 ;
        RECT  1.430 1.930 1.920 2.050 ;
        RECT  1.210 1.930 1.430 2.090 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  0.430 1.930 0.670 2.090 ;
    END
END AOI33D1

MACRO AOI33D2
    CLASS CORE ;
    FOREIGN AOI33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.430 1.370 0.590 ;
        RECT  1.370 0.470 3.385 0.590 ;
        RECT  3.385 0.430 3.605 0.590 ;
        RECT  2.590 1.620 4.570 1.780 ;
        RECT  3.605 0.470 4.570 0.590 ;
        RECT  4.570 0.470 4.710 1.780 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        RECT  0.250 0.725 2.030 0.845 ;
        RECT  2.030 0.725 2.190 1.250 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.750 1.235 ;
        RECT  0.750 1.005 0.870 1.475 ;
        RECT  0.870 1.355 1.680 1.475 ;
        RECT  1.650 0.965 1.680 1.100 ;
        RECT  1.680 0.965 1.840 1.475 ;
        RECT  1.840 0.965 1.870 1.100 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.670 1.235 ;
        RECT  2.670 1.005 2.790 1.475 ;
        RECT  2.790 1.355 4.290 1.475 ;
        RECT  4.290 0.910 4.450 1.475 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 0.930 2.970 1.150 ;
        RECT  2.970 0.725 3.110 1.235 ;
        RECT  3.110 0.725 3.930 0.845 ;
        RECT  3.930 0.725 4.090 1.170 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 2.250 0.300 ;
        RECT  2.250 -0.300 2.470 0.340 ;
        RECT  2.470 -0.300 4.430 0.300 ;
        RECT  4.430 -0.300 4.650 0.340 ;
        RECT  4.650 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 1.920 0.790 2.040 ;
        RECT  0.790 1.620 1.010 2.040 ;
        RECT  1.010 1.920 1.510 2.040 ;
        RECT  1.510 1.620 1.730 2.040 ;
        RECT  1.730 1.920 2.230 2.040 ;
        RECT  2.230 1.620 2.450 2.040 ;
        RECT  2.450 1.920 2.990 2.040 ;
        RECT  2.990 1.900 3.210 2.060 ;
        RECT  3.210 1.900 3.750 2.040 ;
        RECT  3.750 1.900 3.970 2.060 ;
        RECT  3.970 1.900 4.510 2.040 ;
        RECT  4.510 1.900 4.730 2.060 ;
        RECT  0.070 1.620 0.290 2.040 ;
    END
END AOI33D2

MACRO AOI33D4
    CLASS CORE ;
    FOREIGN AOI33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.640 2.830 2.020 ;
        RECT  2.610 0.760 2.830 0.920 ;
        RECT  2.830 0.760 3.250 2.020 ;
        RECT  3.250 1.640 3.630 2.020 ;
        RECT  3.250 0.760 3.630 0.920 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.830 1.270 ;
        RECT  1.830 1.050 1.880 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.530 1.270 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.290 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.725 1.200 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 2.220 0.300 ;
        RECT  2.220 -0.300 2.440 0.340 ;
        RECT  2.440 -0.300 3.020 0.300 ;
        RECT  3.020 -0.300 3.240 0.340 ;
        RECT  3.240 -0.300 3.800 0.300 ;
        RECT  3.800 -0.300 4.020 0.340 ;
        RECT  4.020 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 3.800 2.820 ;
        RECT  3.800 2.180 4.020 2.820 ;
        RECT  4.020 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.405 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.100 1.270 ;
        RECT  0.670 1.930 1.210 2.050 ;
        RECT  1.210 1.930 1.240 2.100 ;
        RECT  1.240 1.390 1.400 2.100 ;
        RECT  1.400 1.930 1.430 2.100 ;
        RECT  1.430 1.930 1.930 2.050 ;
        RECT  1.930 1.930 1.960 2.100 ;
        RECT  1.960 1.370 2.120 2.100 ;
        RECT  2.120 1.960 2.150 2.100 ;
        RECT  1.185 0.430 1.405 0.590 ;
        RECT  0.540 0.470 1.185 0.590 ;
        RECT  0.830 1.410 1.050 1.810 ;
        RECT  0.540 1.410 0.830 1.530 ;
        RECT  0.420 0.470 0.540 1.530 ;
        RECT  0.290 1.410 0.420 1.530 ;
        RECT  4.380 1.960 4.410 2.100 ;
        RECT  4.220 0.420 4.380 2.100 ;
        RECT  3.750 1.390 4.220 1.510 ;
        RECT  4.190 1.960 4.220 2.100 ;
        RECT  3.590 1.050 3.750 1.510 ;
        RECT  0.070 1.410 0.290 1.830 ;
        RECT  0.450 1.670 0.670 2.090 ;
        LAYER M1 ;
        RECT  3.465 1.640 3.630 2.020 ;
        RECT  3.465 0.760 3.630 0.920 ;
    END
END AOI33D4

MACRO BENCD1
    CLASS CORE ;
    FOREIGN BENCD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.940 0.090 2.100 ;
        RECT  0.090 0.420 0.230 2.100 ;
        RECT  0.230 1.390 0.260 2.100 ;
        RECT  0.230 0.420 0.260 0.900 ;
        RECT  0.260 1.940 0.290 2.100 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 0.730 5.030 1.560 ;
        RECT  5.030 1.400 5.190 1.560 ;
        RECT  5.030 0.730 5.280 0.870 ;
        RECT  5.280 0.710 5.520 0.870 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.725 2.970 0.870 ;
        RECT  2.970 0.725 3.110 1.295 ;
        RECT  3.110 1.175 3.330 1.295 ;
        RECT  3.330 1.075 3.470 1.295 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.190 2.020 1.330 ;
        RECT  2.020 1.190 2.330 1.310 ;
        RECT  2.330 1.005 2.470 1.310 ;
        RECT  2.470 1.190 2.620 1.310 ;
        RECT  2.620 1.005 2.790 1.310 ;
        RECT  2.790 1.140 2.840 1.310 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 0.710 3.430 0.955 ;
        RECT  3.470 1.420 3.590 1.560 ;
        RECT  3.430 0.835 3.590 0.955 ;
        RECT  3.590 0.835 3.610 1.560 ;
        RECT  3.610 0.725 3.710 1.560 ;
        RECT  3.710 0.725 3.750 0.955 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 2.050 0.300 ;
        RECT  2.050 -0.300 2.270 0.510 ;
        RECT  2.270 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 2.050 2.820 ;
        RECT  2.050 1.980 2.270 2.820 ;
        RECT  2.270 2.220 2.810 2.820 ;
        RECT  2.810 2.180 3.030 2.820 ;
        RECT  3.030 2.220 3.890 2.820 ;
        RECT  3.890 2.180 4.110 2.820 ;
        RECT  4.110 2.220 5.680 2.820 ;
        RECT  5.680 2.180 5.900 2.820 ;
        RECT  5.900 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.120 0.470 5.660 0.590 ;
        RECT  5.660 0.450 5.880 0.870 ;
        RECT  0.860 1.690 1.680 1.810 ;
        RECT  0.860 0.710 1.680 0.830 ;
        RECT  1.680 0.580 1.820 0.830 ;
        RECT  1.680 1.690 1.840 1.930 ;
        RECT  1.840 1.690 2.600 1.810 ;
        RECT  2.600 1.690 2.720 2.050 ;
        RECT  2.720 1.930 5.570 2.050 ;
        RECT  5.570 1.030 5.730 2.050 ;
        RECT  1.520 0.950 1.640 1.570 ;
        RECT  1.640 0.950 1.940 1.070 ;
        RECT  1.940 0.660 2.060 1.070 ;
        RECT  2.060 0.660 2.390 0.780 ;
        RECT  1.640 1.450 2.450 1.570 ;
        RECT  2.390 0.450 2.510 0.780 ;
        RECT  2.450 1.430 2.680 1.570 ;
        RECT  2.510 0.450 2.680 0.590 ;
        RECT  2.680 1.450 2.840 1.570 ;
        RECT  2.840 1.450 2.960 1.810 ;
        RECT  2.960 1.690 5.310 1.810 ;
        RECT  5.170 1.050 5.310 1.270 ;
        RECT  5.310 1.050 5.430 1.810 ;
        RECT  3.925 0.760 4.045 1.540 ;
        RECT  4.045 0.760 4.260 0.880 ;
        RECT  4.045 1.400 4.280 1.540 ;
        RECT  4.260 0.460 4.480 0.880 ;
        RECT  4.280 1.400 4.520 1.560 ;
        RECT  3.030 0.470 3.570 0.590 ;
        RECT  3.570 0.450 3.810 0.590 ;
        RECT  0.420 0.470 0.540 2.050 ;
        RECT  0.540 0.470 1.250 0.590 ;
        RECT  0.540 1.930 1.260 2.050 ;
        RECT  1.250 0.450 1.490 0.590 ;
        RECT  1.260 1.930 1.500 2.090 ;
        RECT  4.880 0.450 5.120 0.610 ;
        RECT  0.700 0.710 0.860 1.810 ;
        RECT  1.400 1.190 1.520 1.350 ;
        RECT  3.830 1.075 3.925 1.295 ;
        RECT  2.810 0.450 3.030 0.590 ;
        RECT  0.380 1.050 0.420 1.270 ;
    END
END BENCD1

MACRO BENCD2
    CLASS CORE ;
    FOREIGN BENCD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.830 0.230 1.660 ;
        RECT  0.230 1.540 0.450 1.660 ;
        RECT  0.230 0.830 0.460 0.950 ;
        RECT  0.450 1.540 0.610 2.040 ;
        RECT  0.460 0.450 0.620 0.950 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.700 1.380 6.860 1.620 ;
        RECT  6.860 1.380 7.730 1.500 ;
        RECT  7.680 0.710 7.920 0.870 ;
        RECT  7.730 1.380 7.950 1.550 ;
        RECT  7.950 1.380 8.090 1.520 ;
        RECT  7.920 0.730 8.090 0.870 ;
        RECT  8.090 0.730 8.230 1.520 ;
        RECT  8.230 0.730 8.460 0.870 ;
        RECT  8.460 0.710 8.700 0.870 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.670 1.235 ;
        RECT  5.670 1.055 5.850 1.215 ;
        RECT  5.850 1.005 5.990 1.235 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.900 0.720 3.120 0.870 ;
        RECT  3.120 0.750 3.310 0.870 ;
        RECT  3.310 0.750 3.430 1.125 ;
        RECT  3.430 1.005 3.930 1.125 ;
        RECT  3.930 1.005 4.390 1.235 ;
        RECT  4.390 1.075 4.620 1.235 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.190 2.290 1.330 ;
        RECT  2.290 1.190 2.650 1.310 ;
        RECT  2.650 1.005 2.790 1.310 ;
        RECT  2.790 1.140 2.970 1.310 ;
        RECT  2.970 1.005 3.110 1.310 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.550 0.710 3.770 0.870 ;
        RECT  3.770 0.730 4.310 0.850 ;
        RECT  4.310 0.710 4.530 0.870 ;
        RECT  4.530 0.725 4.890 0.850 ;
        RECT  4.890 0.725 4.910 1.350 ;
        RECT  4.910 0.725 5.030 1.560 ;
        RECT  5.030 1.400 5.140 1.560 ;
        RECT  5.140 1.420 5.620 1.540 ;
        RECT  5.620 1.400 5.840 1.560 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.510 ;
        RECT  2.540 -0.300 5.090 0.300 ;
        RECT  5.090 -0.300 5.310 0.340 ;
        RECT  5.310 -0.300 6.920 0.300 ;
        RECT  6.920 -0.300 7.140 0.340 ;
        RECT  7.140 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.350 2.820 ;
        RECT  2.350 1.930 2.510 2.820 ;
        RECT  2.510 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.740 0.470 7.320 0.590 ;
        RECT  7.320 0.450 7.540 0.870 ;
        RECT  7.540 0.470 8.075 0.590 ;
        RECT  8.075 0.470 8.080 0.610 ;
        RECT  8.080 0.450 8.300 0.610 ;
        RECT  8.300 0.470 8.840 0.590 ;
        RECT  8.840 0.470 9.060 0.900 ;
        RECT  7.570 1.930 8.110 2.050 ;
        RECT  8.110 1.910 8.330 2.070 ;
        RECT  8.330 1.930 8.840 2.050 ;
        RECT  8.840 1.630 9.060 2.050 ;
        RECT  1.195 1.690 1.870 1.810 ;
        RECT  1.195 0.710 1.950 0.830 ;
        RECT  1.870 1.690 2.030 1.930 ;
        RECT  1.950 0.580 2.090 0.830 ;
        RECT  2.030 1.690 2.630 1.810 ;
        RECT  2.630 1.690 2.750 2.050 ;
        RECT  2.750 1.930 7.000 2.050 ;
        RECT  7.000 1.670 7.120 2.050 ;
        RECT  7.120 1.670 8.570 1.790 ;
        RECT  8.570 1.030 8.690 1.790 ;
        RECT  8.690 1.030 8.730 1.270 ;
        RECT  1.790 0.950 1.910 1.570 ;
        RECT  1.910 0.950 2.210 1.070 ;
        RECT  2.210 0.660 2.330 1.070 ;
        RECT  2.330 0.660 2.660 0.780 ;
        RECT  1.910 1.450 2.720 1.570 ;
        RECT  2.660 0.450 2.780 0.780 ;
        RECT  2.720 1.430 2.870 1.570 ;
        RECT  2.780 0.450 2.970 0.590 ;
        RECT  2.870 1.430 2.990 1.810 ;
        RECT  2.990 1.690 6.460 1.810 ;
        RECT  6.460 1.080 6.580 1.810 ;
        RECT  6.580 1.080 7.540 1.200 ;
        RECT  7.540 1.040 7.780 1.200 ;
        RECT  5.980 1.400 6.170 1.560 ;
        RECT  5.400 0.750 6.170 0.870 ;
        RECT  6.170 0.450 6.290 1.560 ;
        RECT  6.290 0.450 6.390 0.870 ;
        RECT  3.390 0.470 3.930 0.590 ;
        RECT  3.930 0.450 4.150 0.610 ;
        RECT  4.150 0.470 4.155 0.610 ;
        RECT  4.155 0.470 4.690 0.590 ;
        RECT  4.690 0.450 4.910 0.590 ;
        RECT  4.910 0.470 5.490 0.590 ;
        RECT  5.490 0.450 5.730 0.610 ;
        RECT  3.330 1.450 3.870 1.570 ;
        RECT  3.870 1.430 4.090 1.570 ;
        RECT  4.090 1.450 4.570 1.570 ;
        RECT  4.570 1.430 4.790 1.570 ;
        RECT  0.745 0.470 0.865 2.050 ;
        RECT  0.865 1.930 1.450 2.050 ;
        RECT  0.865 0.470 1.520 0.590 ;
        RECT  1.450 1.930 1.690 2.090 ;
        RECT  1.520 0.450 1.760 0.590 ;
        RECT  7.330 1.910 7.570 2.070 ;
        RECT  1.035 0.710 1.195 1.810 ;
        RECT  1.570 1.190 1.790 1.350 ;
        RECT  5.240 0.750 5.400 1.260 ;
        RECT  3.170 0.450 3.390 0.610 ;
        RECT  3.110 1.430 3.330 1.570 ;
        RECT  0.560 1.080 0.745 1.240 ;
        RECT  6.520 0.450 6.740 0.870 ;
    END
END BENCD2

MACRO BENCD4
    CLASS CORE ;
    FOREIGN BENCD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.650 0.590 2.030 ;
        RECT  0.420 0.490 0.590 0.870 ;
        RECT  0.590 0.490 1.010 2.030 ;
        RECT  1.010 1.650 1.340 2.030 ;
        RECT  1.010 0.490 1.340 0.870 ;
        END
    END X2
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.860 1.380 11.020 1.600 ;
        RECT  11.020 1.380 11.520 1.500 ;
        RECT  11.520 1.380 11.740 1.550 ;
        RECT  11.740 1.380 12.550 1.500 ;
        RECT  12.450 0.710 12.690 0.870 ;
        RECT  12.550 1.380 12.770 1.545 ;
        RECT  12.770 1.380 13.210 1.500 ;
        RECT  12.690 0.730 13.210 0.870 ;
        RECT  13.210 0.730 13.230 1.500 ;
        RECT  13.230 0.710 13.290 1.500 ;
        RECT  13.290 0.710 13.350 1.545 ;
        RECT  13.350 0.710 13.450 0.870 ;
        RECT  13.350 1.380 13.550 1.545 ;
        RECT  13.450 0.730 13.990 0.870 ;
        RECT  13.990 0.710 14.210 0.870 ;
        RECT  14.210 0.730 14.750 0.870 ;
        RECT  14.750 0.710 14.990 0.870 ;
        END
    END S
    PIN M2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.370 1.005 9.510 1.235 ;
        RECT  9.510 1.055 9.690 1.215 ;
        RECT  9.690 1.005 9.830 1.235 ;
        RECT  9.830 1.055 10.030 1.215 ;
        END
    END M2
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.490 0.720 4.730 0.870 ;
        RECT  4.730 0.750 4.920 0.870 ;
        RECT  4.920 0.750 5.040 1.125 ;
        RECT  5.040 1.005 6.490 1.125 ;
        RECT  6.490 1.005 6.950 1.235 ;
        RECT  6.950 1.075 7.145 1.235 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.640 1.190 3.880 1.330 ;
        RECT  3.880 1.190 4.250 1.310 ;
        RECT  4.250 1.005 4.390 1.310 ;
        RECT  4.390 1.140 4.570 1.310 ;
        RECT  4.570 1.005 4.710 1.310 ;
        END
    END M0
    PIN A
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.160 0.710 5.380 0.870 ;
        RECT  5.380 0.730 5.920 0.850 ;
        RECT  5.920 0.710 6.140 0.870 ;
        RECT  6.140 0.730 6.680 0.850 ;
        RECT  6.680 0.710 6.900 0.870 ;
        RECT  6.900 0.730 7.440 0.850 ;
        RECT  7.440 0.710 7.660 0.870 ;
        RECT  8.050 1.400 8.090 1.560 ;
        RECT  7.660 0.730 8.090 0.850 ;
        RECT  8.090 0.730 8.230 1.560 ;
        RECT  8.230 1.400 8.270 1.560 ;
        RECT  8.270 1.420 8.750 1.540 ;
        RECT  8.750 1.400 8.970 1.560 ;
        RECT  8.970 1.420 9.450 1.540 ;
        RECT  9.450 1.400 9.690 1.560 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.160 0.300 ;
        RECT  3.160 -0.300 3.320 0.560 ;
        RECT  3.320 -0.300 3.960 0.300 ;
        RECT  3.960 -0.300 4.120 0.540 ;
        RECT  4.120 -0.300 11.700 0.300 ;
        RECT  11.700 -0.300 11.920 0.340 ;
        RECT  11.920 -0.300 15.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.520 2.820 ;
        RECT  1.520 2.180 1.740 2.820 ;
        RECT  1.740 2.220 3.160 2.820 ;
        RECT  3.160 1.930 3.320 2.820 ;
        RECT  3.320 2.220 3.960 2.820 ;
        RECT  3.960 1.930 4.120 2.820 ;
        RECT  4.120 2.220 5.110 2.820 ;
        RECT  5.110 2.180 5.330 2.820 ;
        RECT  5.330 2.220 5.900 2.820 ;
        RECT  5.900 2.180 6.120 2.820 ;
        RECT  6.120 2.220 15.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  15.130 0.470 15.350 0.895 ;
        RECT  14.590 0.470 15.130 0.590 ;
        RECT  12.390 1.930 12.930 2.050 ;
        RECT  14.370 0.450 14.590 0.610 ;
        RECT  13.830 0.470 14.370 0.590 ;
        RECT  12.930 1.910 13.150 2.070 ;
        RECT  13.150 1.930 13.690 2.050 ;
        RECT  13.610 0.450 13.830 0.610 ;
        RECT  13.690 1.910 13.910 2.070 ;
        RECT  13.910 1.930 14.380 2.050 ;
        RECT  14.380 1.630 14.600 2.050 ;
        RECT  13.070 0.470 13.610 0.590 ;
        RECT  12.850 0.450 13.070 0.610 ;
        RECT  12.310 0.470 12.850 0.590 ;
        RECT  14.600 1.930 15.070 2.050 ;
        RECT  15.070 1.630 15.290 2.050 ;
        RECT  1.860 1.690 2.400 1.810 ;
        RECT  12.090 0.445 12.310 0.865 ;
        RECT  11.530 0.470 12.090 0.590 ;
        RECT  11.310 0.450 11.530 0.870 ;
        RECT  2.400 0.710 2.520 1.810 ;
        RECT  2.520 0.710 2.640 0.830 ;
        RECT  2.520 1.690 2.800 1.810 ;
        RECT  2.640 0.420 2.860 0.830 ;
        RECT  2.800 1.690 2.960 1.930 ;
        RECT  2.960 1.690 3.560 1.810 ;
        RECT  2.860 0.710 3.560 0.830 ;
        RECT  3.560 0.580 3.700 0.830 ;
        RECT  3.560 1.690 3.720 1.930 ;
        RECT  3.720 1.690 4.240 1.810 ;
        RECT  4.240 1.690 4.360 2.050 ;
        RECT  4.360 1.930 11.120 2.050 ;
        RECT  11.120 1.670 11.240 2.050 ;
        RECT  11.240 1.670 13.920 1.790 ;
        RECT  13.920 1.080 14.040 1.790 ;
        RECT  14.040 1.080 14.700 1.240 ;
        RECT  2.780 0.950 2.940 1.570 ;
        RECT  2.940 0.950 3.820 1.070 ;
        RECT  3.820 0.660 3.940 1.070 ;
        RECT  3.940 0.660 4.240 0.780 ;
        RECT  2.940 1.450 4.330 1.570 ;
        RECT  4.240 0.450 4.360 0.780 ;
        RECT  4.330 1.430 4.480 1.570 ;
        RECT  4.360 0.450 4.570 0.590 ;
        RECT  4.480 1.430 4.600 1.810 ;
        RECT  4.600 1.690 10.620 1.810 ;
        RECT  10.620 1.080 10.740 1.810 ;
        RECT  10.740 1.080 12.860 1.240 ;
        RECT  9.050 0.750 9.170 1.210 ;
        RECT  9.170 0.750 9.920 0.870 ;
        RECT  9.920 0.450 10.140 0.870 ;
        RECT  10.120 1.400 10.240 1.560 ;
        RECT  10.140 0.750 10.240 0.870 ;
        RECT  10.240 0.750 10.360 1.560 ;
        RECT  5.000 0.470 5.540 0.590 ;
        RECT  5.540 0.450 5.760 0.610 ;
        RECT  5.760 0.470 5.765 0.610 ;
        RECT  5.765 0.470 6.300 0.590 ;
        RECT  6.300 0.450 6.520 0.610 ;
        RECT  6.520 0.470 7.060 0.590 ;
        RECT  7.060 0.450 7.280 0.610 ;
        RECT  7.280 0.470 7.820 0.590 ;
        RECT  7.820 0.450 8.040 0.610 ;
        RECT  8.040 0.470 8.520 0.590 ;
        RECT  8.520 0.450 8.740 0.610 ;
        RECT  8.740 0.470 9.220 0.590 ;
        RECT  9.220 0.450 9.460 0.610 ;
        RECT  4.940 1.450 5.500 1.570 ;
        RECT  5.500 1.410 5.720 1.570 ;
        RECT  5.720 1.450 6.300 1.570 ;
        RECT  6.300 1.410 6.520 1.570 ;
        RECT  6.520 1.450 7.000 1.570 ;
        RECT  7.000 1.410 7.220 1.570 ;
        RECT  7.220 1.450 7.700 1.570 ;
        RECT  7.700 1.410 7.920 1.570 ;
        RECT  1.460 0.470 1.580 2.050 ;
        RECT  1.580 0.470 2.260 0.590 ;
        RECT  1.580 1.930 2.380 2.050 ;
        RECT  2.260 0.450 2.500 0.590 ;
        RECT  2.380 1.930 2.620 2.090 ;
        RECT  1.980 0.710 2.100 1.540 ;
        RECT  2.100 1.400 2.220 1.540 ;
        RECT  10.840 0.470 11.310 0.590 ;
        RECT  12.150 1.910 12.390 2.070 ;
        RECT  1.710 1.030 1.860 1.810 ;
        RECT  8.670 1.050 9.050 1.210 ;
        RECT  4.780 0.450 5.000 0.610 ;
        RECT  4.720 1.430 4.940 1.570 ;
        RECT  1.250 1.080 1.460 1.240 ;
        RECT  1.860 0.710 1.980 0.870 ;
        RECT  10.620 0.450 10.840 0.870 ;
        LAYER M1 ;
        RECT  1.225 0.490 1.340 0.870 ;
        RECT  1.225 1.650 1.340 2.030 ;
    END
END BENCD4

MACRO BHD
    CLASS CORE ;
    FOREIGN BHD 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION INOUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.040 0.420 1.280 ;
        RECT  0.420 1.040 0.470 1.930 ;
        RECT  0.470 1.160 0.540 1.930 ;
        RECT  0.540 1.810 1.020 1.930 ;
        RECT  1.020 0.570 1.190 1.930 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.210 1.390 0.250 2.050 ;
        RECT  0.210 0.520 0.250 0.920 ;
        RECT  0.250 0.800 0.710 0.920 ;
        RECT  0.710 0.800 0.870 1.290 ;
        RECT  0.090 0.520 0.210 2.050 ;
    END
END BHD

MACRO BMLD1
    CLASS CORE ;
    FOREIGN BMLD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.445 0.550 0.990 ;
        RECT  0.550 0.865 0.610 0.990 ;
        RECT  0.610 0.865 0.770 1.270 ;
        END
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.230 0.725 4.390 1.285 ;
        END
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.060 0.835 0.090 1.685 ;
        RECT  0.090 0.420 0.180 2.070 ;
        RECT  0.180 1.565 0.250 2.070 ;
        RECT  0.180 0.420 0.250 0.955 ;
        END
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.950 0.865 6.110 1.270 ;
        RECT  6.110 0.865 6.170 0.990 ;
        RECT  6.170 0.445 6.310 0.990 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.445 2.410 0.990 ;
        RECT  2.410 0.445 2.470 1.270 ;
        RECT  2.470 0.865 2.570 1.270 ;
        END
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.005 4.070 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.060 1.930 1.300 2.070 ;
        RECT  2.110 1.090 2.200 1.520 ;
        RECT  2.940 1.350 3.040 1.570 ;
        RECT  3.620 0.720 3.750 1.810 ;
        RECT  5.610 1.000 5.700 1.220 ;
        RECT  4.990 0.710 5.130 1.810 ;
        RECT  1.300 1.930 6.470 2.050 ;
        RECT  6.470 1.570 6.540 2.050 ;
        RECT  6.470 0.420 6.540 0.915 ;
        RECT  6.540 0.420 6.660 2.050 ;
        RECT  5.130 1.690 6.230 1.810 ;
        RECT  6.230 1.110 6.350 1.810 ;
        RECT  6.350 1.110 6.420 1.330 ;
        RECT  5.700 0.565 5.820 1.570 ;
        RECT  5.820 1.410 5.940 1.570 ;
        RECT  5.820 0.565 5.940 0.725 ;
        RECT  3.750 1.670 3.880 1.810 ;
        RECT  3.750 0.720 3.920 0.880 ;
        RECT  3.880 1.690 4.750 1.810 ;
        RECT  4.750 0.470 4.870 1.810 ;
        RECT  4.870 0.470 5.330 0.590 ;
        RECT  5.330 0.470 5.460 1.570 ;
        RECT  5.460 1.400 5.570 1.570 ;
        RECT  5.460 0.470 5.570 0.630 ;
        RECT  2.940 0.610 3.040 0.830 ;
        RECT  3.040 0.470 3.160 1.570 ;
        RECT  4.390 1.410 4.510 1.570 ;
        RECT  3.160 0.470 4.510 0.590 ;
        RECT  4.510 0.470 4.630 1.570 ;
        RECT  2.200 1.090 2.250 1.810 ;
        RECT  2.250 1.400 2.320 1.810 ;
        RECT  2.320 1.690 3.280 1.810 ;
        RECT  3.280 1.670 3.360 1.810 ;
        RECT  3.280 0.720 3.360 0.880 ;
        RECT  3.360 0.720 3.500 1.810 ;
        RECT  2.590 0.470 2.700 0.690 ;
        RECT  2.700 0.470 2.820 1.570 ;
        RECT  2.820 1.035 2.920 1.195 ;
        RECT  1.980 0.440 2.050 0.955 ;
        RECT  1.980 1.670 2.080 1.810 ;
        RECT  0.370 1.110 0.490 1.810 ;
        RECT  0.490 1.690 1.480 1.810 ;
        RECT  1.480 1.670 1.600 1.810 ;
        RECT  1.500 0.610 1.600 0.830 ;
        RECT  1.600 0.610 1.740 1.810 ;
        RECT  1.140 0.610 1.240 0.830 ;
        RECT  1.240 0.610 1.360 1.570 ;
        RECT  0.730 0.550 0.900 0.710 ;
        RECT  0.900 0.550 1.020 1.570 ;
        RECT  1.020 1.035 1.120 1.195 ;
        RECT  2.530 1.410 2.700 1.570 ;
        RECT  1.860 0.440 1.980 1.810 ;
        RECT  0.310 1.110 0.370 1.330 ;
        RECT  1.140 1.350 1.240 1.570 ;
        RECT  0.730 1.410 0.900 1.570 ;
    END
END BMLD1

MACRO BMLD2
    CLASS CORE ;
    FOREIGN BMLD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.445 1.190 0.990 ;
        RECT  1.190 0.865 1.250 0.990 ;
        RECT  1.250 0.865 1.410 1.270 ;
        END
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.870 0.725 5.030 1.285 ;
        END
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.835 0.550 1.685 ;
        RECT  0.550 1.565 0.590 1.685 ;
        RECT  0.550 0.835 0.590 0.955 ;
        RECT  0.590 1.565 0.750 2.070 ;
        RECT  0.590 0.420 0.750 0.955 ;
        END
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.590 0.830 6.750 1.270 ;
        RECT  6.750 0.830 6.810 0.955 ;
        RECT  6.810 0.445 6.950 0.955 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.445 3.050 0.955 ;
        RECT  3.050 0.445 3.110 1.270 ;
        RECT  3.110 0.830 3.210 1.270 ;
        END
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.005 4.710 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 0.970 0.300 ;
        RECT  0.970 -0.300 1.190 0.325 ;
        RECT  1.190 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 0.970 2.820 ;
        RECT  0.970 2.180 1.190 2.820 ;
        RECT  1.190 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 1.930 7.110 2.050 ;
        RECT  7.110 1.570 7.180 2.050 ;
        RECT  7.110 0.420 7.180 0.915 ;
        RECT  7.180 0.420 7.300 2.050 ;
        RECT  5.770 1.690 6.870 1.810 ;
        RECT  6.870 1.110 6.990 1.810 ;
        RECT  6.990 1.110 7.060 1.330 ;
        RECT  6.340 0.460 6.460 1.570 ;
        RECT  6.460 1.410 6.580 1.570 ;
        RECT  6.460 0.460 6.580 0.620 ;
        RECT  4.390 1.665 4.520 1.810 ;
        RECT  4.390 0.720 4.560 0.880 ;
        RECT  4.520 1.690 5.390 1.810 ;
        RECT  5.390 0.470 5.510 1.810 ;
        RECT  5.510 0.470 5.970 0.590 ;
        RECT  5.970 0.470 6.100 1.570 ;
        RECT  6.100 1.410 6.210 1.570 ;
        RECT  6.100 0.470 6.210 0.630 ;
        RECT  3.580 0.610 3.680 0.830 ;
        RECT  3.680 0.470 3.800 1.570 ;
        RECT  5.030 1.410 5.150 1.570 ;
        RECT  3.800 0.470 5.150 0.590 ;
        RECT  5.150 0.470 5.270 1.570 ;
        RECT  2.840 1.090 2.890 1.810 ;
        RECT  2.890 1.400 2.960 1.810 ;
        RECT  2.960 1.690 3.920 1.810 ;
        RECT  3.920 1.670 4.000 1.810 ;
        RECT  3.920 0.720 4.000 0.880 ;
        RECT  4.000 0.720 4.140 1.810 ;
        RECT  3.230 0.470 3.340 0.690 ;
        RECT  3.340 0.470 3.460 1.570 ;
        RECT  3.460 1.035 3.560 1.195 ;
        RECT  2.620 0.440 2.690 0.955 ;
        RECT  2.620 1.670 2.720 1.810 ;
        RECT  1.010 1.140 1.130 1.810 ;
        RECT  1.130 1.690 2.120 1.810 ;
        RECT  2.120 1.670 2.240 1.810 ;
        RECT  2.140 0.610 2.240 0.830 ;
        RECT  2.240 0.610 2.380 1.810 ;
        RECT  1.780 0.610 1.880 0.830 ;
        RECT  1.880 0.610 2.000 1.570 ;
        RECT  1.370 0.550 1.540 0.710 ;
        RECT  1.540 0.550 1.660 1.570 ;
        RECT  1.660 1.035 1.760 1.195 ;
        RECT  5.630 0.710 5.770 1.810 ;
        RECT  6.250 1.000 6.340 1.220 ;
        RECT  4.260 0.720 4.390 1.810 ;
        RECT  3.580 1.350 3.680 1.570 ;
        RECT  2.750 1.090 2.840 1.520 ;
        RECT  1.700 1.930 1.940 2.070 ;
        RECT  3.170 1.410 3.340 1.570 ;
        RECT  2.500 0.440 2.620 1.810 ;
        RECT  0.690 1.140 1.010 1.300 ;
        RECT  1.780 1.350 1.880 1.570 ;
        RECT  1.370 1.410 1.540 1.570 ;
    END
END BMLD2

MACRO BMLD4
    CLASS CORE ;
    FOREIGN BMLD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN X2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.290 0.830 8.410 1.270 ;
        RECT  8.410 0.445 8.450 1.270 ;
        RECT  8.450 0.445 8.550 0.955 ;
        END
    END X2
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END S
    PIN PP
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.810 1.650 9.230 2.030 ;
        RECT  8.810 0.490 9.230 0.870 ;
        RECT  9.230 0.490 9.650 2.030 ;
        RECT  9.650 1.650 9.780 2.030 ;
        RECT  9.650 0.490 9.780 0.870 ;
        END
    END PP
    PIN M1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.445 0.870 0.955 ;
        RECT  0.870 0.830 0.970 0.955 ;
        RECT  0.970 0.830 1.130 1.290 ;
        END
    END M1
    PIN M0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.810 1.005 6.310 1.235 ;
        END
    END M0
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.420 0.300 ;
        RECT  8.420 -0.300 8.640 0.320 ;
        RECT  8.640 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.420 2.820 ;
        RECT  8.420 2.180 8.640 2.820 ;
        RECT  8.640 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.800 0.720 4.580 0.880 ;
        RECT  4.580 0.720 4.710 1.810 ;
        RECT  0.730 1.075 0.850 1.810 ;
        RECT  0.850 1.690 1.950 1.810 ;
        RECT  1.950 0.710 2.090 1.810 ;
        RECT  1.140 0.470 1.260 0.630 ;
        RECT  1.260 0.470 1.380 1.570 ;
        RECT  1.380 1.045 1.470 1.265 ;
        RECT  3.840 1.665 4.580 1.810 ;
        RECT  2.330 1.690 3.840 1.810 ;
        RECT  2.210 0.470 2.330 1.810 ;
        RECT  1.750 0.470 2.210 0.590 ;
        RECT  1.620 0.470 1.750 1.570 ;
        RECT  1.510 0.470 1.620 0.630 ;
        RECT  5.320 0.610 5.440 0.830 ;
        RECT  5.320 1.350 5.440 1.570 ;
        RECT  5.200 0.470 5.320 1.570 ;
        RECT  3.310 0.470 5.200 0.590 ;
        RECT  2.570 1.410 3.380 1.570 ;
        RECT  2.570 0.470 3.310 0.630 ;
        RECT  5.680 1.410 5.830 1.570 ;
        RECT  5.680 0.420 5.810 0.840 ;
        RECT  5.590 0.420 5.680 1.570 ;
        RECT  5.560 0.720 5.590 1.570 ;
        RECT  6.440 1.030 6.600 1.480 ;
        RECT  6.160 1.360 6.440 1.480 ;
        RECT  6.040 1.360 6.160 1.810 ;
        RECT  5.080 1.690 6.040 1.810 ;
        RECT  5.000 0.720 5.080 0.880 ;
        RECT  5.000 1.670 5.080 1.810 ;
        RECT  7.020 0.550 7.140 1.810 ;
        RECT  6.500 0.550 7.020 0.710 ;
        RECT  6.280 1.650 7.020 1.810 ;
        RECT  7.810 0.640 7.910 0.800 ;
        RECT  7.810 1.410 7.910 1.570 ;
        RECT  7.680 1.930 7.920 2.070 ;
        RECT  0.610 1.930 7.680 2.050 ;
        RECT  0.530 0.420 0.610 0.920 ;
        RECT  0.530 1.570 0.610 2.050 ;
        RECT  0.450 0.420 0.530 2.050 ;
        RECT  8.150 0.550 8.270 0.710 ;
        RECT  8.150 1.410 8.270 1.570 ;
        RECT  8.030 0.550 8.150 1.570 ;
        RECT  8.690 1.080 8.900 1.240 ;
        RECT  8.570 1.080 8.690 1.810 ;
        RECT  7.520 1.690 8.570 1.810 ;
        RECT  7.400 0.640 7.550 0.800 ;
        RECT  7.400 1.670 7.520 1.810 ;
        RECT  7.930 1.035 8.030 1.195 ;
        RECT  0.410 0.800 0.450 1.690 ;
        RECT  7.690 0.640 7.810 1.570 ;
        RECT  6.280 0.420 6.500 0.840 ;
        RECT  4.860 0.720 5.000 1.810 ;
        RECT  5.440 1.035 5.560 1.195 ;
        RECT  2.450 0.470 2.570 1.570 ;
        RECT  1.510 1.410 1.620 1.570 ;
        RECT  0.650 1.075 0.730 1.295 ;
        RECT  7.260 0.640 7.400 1.810 ;
        RECT  1.140 1.410 1.260 1.570 ;
        LAYER M1 ;
        RECT  8.810 1.650 9.015 2.030 ;
        RECT  8.810 0.490 9.015 0.870 ;
    END
END BMLD4

MACRO BUFFD0
    CLASS CORE ;
    FOREIGN BUFFD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.420 0.600 0.590 ;
        RECT  0.360 1.915 0.730 2.075 ;
        RECT  0.600 0.470 0.730 0.590 ;
        RECT  0.730 1.565 0.740 2.075 ;
        RECT  0.730 0.470 0.740 0.955 ;
        RECT  0.740 0.470 0.870 2.075 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.550 1.050 0.620 1.270 ;
        RECT  0.390 0.710 0.550 1.635 ;
    END
END BUFFD0

MACRO BUFFD1
    CLASS CORE ;
    FOREIGN BUFFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.960 1.030 2.100 ;
        RECT  1.030 0.420 1.190 2.100 ;
        RECT  1.190 1.960 1.220 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.340 ;
        RECT  0.760 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 2.180 0.760 2.820 ;
        RECT  0.760 2.220 1.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.720 0.470 0.880 2.050 ;
        RECT  0.100 0.470 0.720 0.630 ;
        RECT  0.100 1.890 0.720 2.050 ;
    END
END BUFFD1

MACRO BUFFD12
    CLASS CORE ;
    FOREIGN BUFFD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.640 3.150 2.020 ;
        RECT  1.490 0.500 3.150 0.880 ;
        RECT  3.150 0.500 3.570 2.020 ;
        RECT  3.570 1.640 5.310 2.020 ;
        RECT  3.570 0.500 5.310 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.960 1.080 2.555 1.240 ;
        RECT  0.960 1.960 0.990 2.100 ;
        RECT  0.800 0.420 0.960 2.100 ;
        RECT  0.300 0.750 0.800 0.870 ;
        RECT  0.270 1.650 0.800 1.770 ;
        RECT  0.770 1.960 0.800 2.100 ;
        RECT  0.080 0.450 0.300 0.870 ;
        RECT  0.270 1.960 0.300 2.100 ;
        RECT  0.110 1.370 0.270 2.100 ;
        RECT  0.080 1.960 0.110 2.100 ;
        LAYER M1 ;
        RECT  1.490 0.500 2.935 0.880 ;
        RECT  1.490 1.640 2.935 2.020 ;
        RECT  3.785 0.500 5.310 0.880 ;
        RECT  3.785 1.640 5.310 2.020 ;
    END
END BUFFD12

MACRO BUFFD16
    CLASS CORE ;
    FOREIGN BUFFD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.640 4.110 2.020 ;
        RECT  1.800 0.500 4.110 0.880 ;
        RECT  4.110 0.500 4.530 2.020 ;
        RECT  4.530 1.640 6.930 2.020 ;
        RECT  4.530 0.500 6.930 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.300 1.080 3.220 1.240 ;
        RECT  1.300 1.960 1.330 2.100 ;
        RECT  1.140 0.420 1.300 2.100 ;
        RECT  0.640 0.750 1.140 0.870 ;
        RECT  0.610 1.650 1.140 1.770 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  0.420 0.450 0.640 0.870 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 1.370 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  1.800 0.500 3.895 0.880 ;
        RECT  1.800 1.640 3.895 2.020 ;
        RECT  4.745 0.500 6.930 0.880 ;
        RECT  4.745 1.640 6.930 2.020 ;
    END
END BUFFD16

MACRO BUFFD2
    CLASS CORE ;
    FOREIGN BUFFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.960 0.890 2.100 ;
        RECT  0.890 1.390 1.050 2.100 ;
        RECT  0.890 0.420 1.050 0.900 ;
        RECT  1.050 1.960 1.080 2.100 ;
        RECT  1.050 0.780 1.190 1.515 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.070 1.635 0.290 2.055 ;
        RECT  0.070 0.465 0.290 0.885 ;
        RECT  0.290 1.635 0.610 1.755 ;
        RECT  0.290 0.765 0.610 0.885 ;
        RECT  0.610 0.765 0.770 1.755 ;
    END
END BUFFD2

MACRO BUFFD20
    CLASS CORE ;
    FOREIGN BUFFD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.640 5.390 2.020 ;
        RECT  2.140 0.500 5.390 0.880 ;
        RECT  5.390 0.500 5.810 2.020 ;
        RECT  5.810 1.640 8.840 2.020 ;
        RECT  5.810 0.500 8.840 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.640 1.080 4.030 1.240 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.480 0.420 1.640 2.100 ;
        RECT  0.980 0.750 1.480 0.870 ;
        RECT  0.950 1.635 1.480 1.755 ;
        RECT  1.450 1.960 1.480 2.100 ;
        RECT  0.760 0.450 0.980 0.870 ;
        RECT  0.950 1.960 0.980 2.100 ;
        RECT  0.790 1.370 0.950 2.100 ;
        RECT  0.260 1.635 0.790 1.755 ;
        RECT  0.760 1.960 0.790 2.100 ;
        RECT  0.290 0.750 0.760 0.870 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  2.140 0.500 5.175 0.880 ;
        RECT  2.140 1.640 5.175 2.020 ;
        RECT  6.025 0.500 8.840 0.880 ;
        RECT  6.025 1.640 8.840 2.020 ;
    END
END BUFFD20

MACRO BUFFD24
    CLASS CORE ;
    FOREIGN BUFFD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.640 6.030 2.020 ;
        RECT  2.490 0.500 6.030 0.880 ;
        RECT  6.030 0.500 6.450 2.020 ;
        RECT  6.450 1.640 10.440 2.020 ;
        RECT  6.450 0.500 10.440 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.990 1.080 5.315 1.240 ;
        RECT  1.990 1.960 2.020 2.100 ;
        RECT  1.830 0.420 1.990 2.100 ;
        RECT  1.330 0.750 1.830 0.870 ;
        RECT  1.300 1.650 1.830 1.770 ;
        RECT  1.800 1.960 1.830 2.100 ;
        RECT  1.110 0.450 1.330 0.870 ;
        RECT  1.300 1.960 1.330 2.100 ;
        RECT  1.140 1.370 1.300 2.100 ;
        RECT  0.610 1.650 1.140 1.770 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  0.640 0.750 1.110 0.870 ;
        RECT  0.420 0.450 0.640 0.870 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 1.370 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  2.490 0.500 5.815 0.880 ;
        RECT  2.490 1.640 5.815 2.020 ;
        RECT  6.665 0.500 10.440 0.880 ;
        RECT  6.665 1.640 10.440 2.020 ;
    END
END BUFFD24

MACRO BUFFD3
    CLASS CORE ;
    FOREIGN BUFFD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.640 1.230 2.020 ;
        RECT  0.840 0.500 1.230 0.880 ;
        RECT  1.230 0.500 1.650 2.020 ;
        RECT  1.650 1.640 1.850 2.020 ;
        RECT  1.650 0.500 1.850 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 1.240 0.300 ;
        RECT  1.240 -0.300 1.460 0.340 ;
        RECT  1.460 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.180 0.670 2.820 ;
        RECT  0.670 2.220 1.240 2.820 ;
        RECT  1.240 2.180 1.460 2.820 ;
        RECT  1.460 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.280 0.765 0.400 0.885 ;
        RECT  0.400 0.765 0.520 1.755 ;
        RECT  0.520 1.080 0.950 1.240 ;
        RECT  0.280 1.635 0.400 1.755 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  0.060 1.635 0.280 2.055 ;
        LAYER M1 ;
        RECT  0.840 1.640 1.015 2.020 ;
        RECT  0.840 0.500 1.015 0.880 ;
    END
END BUFFD3

MACRO BUFFD4
    CLASS CORE ;
    FOREIGN BUFFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.650 1.550 2.030 ;
        RECT  1.170 0.490 1.550 0.870 ;
        RECT  1.550 0.490 1.970 2.030 ;
        RECT  1.970 1.650 2.110 2.030 ;
        RECT  1.970 0.490 2.110 0.870 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.640 1.080 1.280 1.240 ;
        RECT  0.640 1.960 0.670 2.100 ;
        RECT  0.480 0.420 0.640 2.100 ;
        RECT  0.450 1.960 0.480 2.100 ;
        LAYER M1 ;
        RECT  1.170 0.490 1.335 0.870 ;
        RECT  1.170 1.650 1.335 2.030 ;
    END
END BUFFD4

MACRO BUFFD6
    CLASS CORE ;
    FOREIGN BUFFD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.640 1.870 2.020 ;
        RECT  1.140 0.500 1.870 0.880 ;
        RECT  1.870 0.500 2.290 2.020 ;
        RECT  2.290 1.640 2.770 2.020 ;
        RECT  2.290 0.500 2.770 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.460 0.420 0.620 2.100 ;
        RECT  0.620 1.960 0.650 2.100 ;
        RECT  0.620 1.080 1.510 1.240 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  2.505 1.640 2.770 2.020 ;
        RECT  2.505 0.500 2.770 0.880 ;
        RECT  1.140 1.640 1.655 2.020 ;
        RECT  1.140 0.500 1.655 0.880 ;
    END
END BUFFD6

MACRO BUFFD8
    CLASS CORE ;
    FOREIGN BUFFD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.640 1.870 2.020 ;
        RECT  1.120 0.500 1.870 0.880 ;
        RECT  1.870 0.500 2.290 2.020 ;
        RECT  2.290 1.640 3.410 2.020 ;
        RECT  2.290 0.500 3.410 0.880 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.620 1.080 1.490 1.240 ;
        RECT  0.620 1.960 0.650 2.100 ;
        RECT  0.460 0.420 0.620 2.100 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  1.120 0.500 1.655 0.880 ;
        RECT  1.120 1.640 1.655 2.020 ;
        RECT  2.505 0.500 3.410 0.880 ;
        RECT  2.505 1.640 3.410 2.020 ;
    END
END BUFFD8

MACRO BUFTD0
    CLASS CORE ;
    FOREIGN BUFTD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.420 2.790 1.950 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.110 0.410 1.330 ;
        RECT  0.410 1.110 0.550 1.515 ;
        RECT  0.550 1.285 0.750 1.515 ;
        RECT  0.750 1.285 0.870 1.930 ;
        RECT  0.870 1.810 1.480 1.930 ;
        RECT  1.480 1.400 1.600 1.930 ;
        RECT  1.600 1.400 1.800 1.520 ;
        RECT  1.800 1.000 1.960 1.520 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.255 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.170 0.300 ;
        RECT  1.170 -0.300 1.390 0.340 ;
        RECT  1.390 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.370 2.820 ;
        RECT  1.370 2.180 1.590 2.820 ;
        RECT  1.590 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.470 2.350 0.590 ;
        RECT  2.350 0.470 2.510 1.010 ;
        RECT  1.800 0.710 2.110 0.870 ;
        RECT  2.110 0.710 2.230 1.900 ;
        RECT  2.230 1.300 2.510 1.460 ;
        RECT  0.210 1.470 0.250 1.710 ;
        RECT  0.210 0.420 0.250 0.960 ;
        RECT  0.250 0.800 0.790 0.960 ;
        RECT  1.050 0.470 1.210 1.690 ;
        RECT  0.750 0.470 1.050 0.630 ;
        RECT  1.750 1.740 2.110 1.900 ;
        RECT  0.090 0.420 0.210 1.710 ;
    END
END BUFTD0

MACRO BUFTD1
    CLASS CORE ;
    FOREIGN BUFTD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.465 2.790 2.070 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.110 0.410 1.330 ;
        RECT  0.410 1.110 0.550 1.515 ;
        RECT  0.550 1.285 0.710 1.515 ;
        RECT  0.710 1.285 0.850 2.050 ;
        RECT  0.850 1.285 0.870 1.515 ;
        RECT  0.850 1.930 1.480 2.050 ;
        RECT  1.480 1.455 1.600 2.050 ;
        RECT  1.600 1.455 1.800 1.575 ;
        RECT  1.800 1.000 1.960 1.575 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.255 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.170 0.300 ;
        RECT  1.170 -0.300 1.390 0.340 ;
        RECT  1.390 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 1.370 2.820 ;
        RECT  1.370 2.180 1.590 2.820 ;
        RECT  1.590 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.995 0.470 1.020 0.590 ;
        RECT  1.020 0.470 1.140 1.810 ;
        RECT  1.140 1.410 1.240 1.810 ;
        RECT  1.140 0.470 2.350 0.590 ;
        RECT  2.350 0.470 2.510 1.110 ;
        RECT  1.800 0.710 2.110 0.870 ;
        RECT  2.110 0.710 2.230 2.020 ;
        RECT  2.230 1.240 2.510 1.400 ;
        RECT  0.210 1.470 0.250 1.710 ;
        RECT  0.210 0.420 0.250 0.960 ;
        RECT  0.250 0.800 0.790 0.960 ;
        RECT  0.750 0.430 0.995 0.590 ;
        RECT  1.750 1.860 2.110 2.020 ;
        RECT  0.090 0.420 0.210 1.710 ;
    END
END BUFTD1

MACRO BUFTD12
    CLASS CORE ;
    FOREIGN BUFTD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.640 5.070 2.020 ;
        RECT  3.400 0.480 5.070 0.640 ;
        RECT  5.070 0.480 5.490 2.020 ;
        RECT  5.490 1.640 7.240 2.020 ;
        RECT  5.490 0.480 7.260 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.030 0.490 2.050 ;
        RECT  0.490 1.930 1.700 2.050 ;
        RECT  1.700 1.395 1.820 2.050 ;
        RECT  1.820 1.395 2.330 1.515 ;
        RECT  2.330 1.005 2.450 1.515 ;
        RECT  2.450 1.005 2.790 1.235 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.880 1.510 1.810 ;
        RECT  1.105 0.880 1.390 1.040 ;
        RECT  0.745 1.690 1.390 1.810 ;
        RECT  0.625 0.790 0.745 1.810 ;
        RECT  0.250 0.790 0.625 0.910 ;
        RECT  0.230 0.430 0.250 0.910 ;
        RECT  3.290 1.170 3.530 1.330 ;
        RECT  3.030 1.190 3.290 1.330 ;
        RECT  2.910 0.710 3.030 1.510 ;
        RECT  2.890 1.960 2.920 2.100 ;
        RECT  2.395 0.710 2.910 0.870 ;
        RECT  2.890 1.390 2.910 1.510 ;
        RECT  2.730 1.390 2.890 2.100 ;
        RECT  2.700 1.930 2.730 2.100 ;
        RECT  2.220 1.930 2.700 2.050 ;
        RECT  2.190 1.930 2.220 2.090 ;
        RECT  2.030 1.640 2.190 2.090 ;
        RECT  3.650 0.930 3.890 1.090 ;
        RECT  3.270 0.930 3.650 1.050 ;
        RECT  3.150 0.470 3.270 1.050 ;
        RECT  1.680 0.470 3.150 0.590 ;
        RECT  1.460 0.430 1.680 0.590 ;
        RECT  0.990 0.470 1.460 0.590 ;
        RECT  0.985 1.410 1.260 1.570 ;
        RECT  0.985 0.430 0.990 0.590 ;
        RECT  0.865 0.430 0.985 1.570 ;
        RECT  0.750 0.430 0.865 0.590 ;
        RECT  2.000 1.930 2.030 2.090 ;
        RECT  0.090 0.430 0.230 1.690 ;
        LAYER M1 ;
        RECT  3.400 0.480 4.855 0.640 ;
        RECT  3.420 1.640 4.855 2.020 ;
        RECT  5.705 0.480 7.260 0.640 ;
        RECT  5.705 1.640 7.240 2.020 ;
    END
END BUFTD12

MACRO BUFTD16
    CLASS CORE ;
    FOREIGN BUFTD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.410 1.640 5.710 2.020 ;
        RECT  3.390 0.480 5.710 0.640 ;
        RECT  5.710 0.480 6.130 2.020 ;
        RECT  6.130 1.640 8.530 2.020 ;
        RECT  6.130 0.480 8.550 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.030 0.490 2.050 ;
        RECT  0.490 1.930 1.700 2.050 ;
        RECT  1.700 1.395 1.820 2.050 ;
        RECT  1.820 1.395 2.330 1.515 ;
        RECT  2.330 1.005 2.450 1.515 ;
        RECT  2.450 1.005 2.790 1.235 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.880 1.510 1.810 ;
        RECT  1.105 0.880 1.390 1.040 ;
        RECT  0.745 1.690 1.390 1.810 ;
        RECT  0.625 0.790 0.745 1.810 ;
        RECT  0.250 0.790 0.625 0.910 ;
        RECT  0.230 0.485 0.250 0.910 ;
        RECT  3.280 1.180 3.520 1.330 ;
        RECT  3.030 1.210 3.280 1.330 ;
        RECT  2.910 0.710 3.030 1.510 ;
        RECT  2.890 1.960 2.920 2.100 ;
        RECT  2.395 0.710 2.910 0.870 ;
        RECT  2.890 1.390 2.910 1.510 ;
        RECT  2.730 1.390 2.890 2.100 ;
        RECT  2.700 1.930 2.730 2.100 ;
        RECT  2.220 1.930 2.700 2.050 ;
        RECT  2.190 1.930 2.220 2.090 ;
        RECT  2.030 1.640 2.190 2.090 ;
        RECT  3.980 0.940 4.220 1.100 ;
        RECT  3.270 0.940 3.980 1.060 ;
        RECT  3.150 0.470 3.270 1.060 ;
        RECT  1.680 0.470 3.150 0.590 ;
        RECT  1.460 0.430 1.680 0.590 ;
        RECT  0.990 0.470 1.460 0.590 ;
        RECT  0.985 1.410 1.260 1.570 ;
        RECT  0.985 0.430 0.990 0.590 ;
        RECT  0.865 0.430 0.985 1.570 ;
        RECT  0.750 0.430 0.865 0.590 ;
        RECT  2.000 1.930 2.030 2.090 ;
        RECT  0.090 0.485 0.230 2.040 ;
        LAYER M1 ;
        RECT  3.390 0.480 5.495 0.640 ;
        RECT  3.410 1.640 5.495 2.020 ;
        RECT  6.345 0.480 8.550 0.640 ;
        RECT  6.345 1.640 8.530 2.020 ;
    END
END BUFTD16

MACRO BUFTD2
    CLASS CORE ;
    FOREIGN BUFTD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.555 2.690 2.055 ;
        RECT  2.690 1.555 2.970 1.675 ;
        RECT  2.500 0.520 2.970 0.680 ;
        RECT  2.970 0.520 3.110 1.675 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.110 0.410 1.330 ;
        RECT  0.410 1.110 0.550 1.515 ;
        RECT  0.550 1.285 0.710 1.515 ;
        RECT  0.710 1.285 0.850 2.050 ;
        RECT  0.850 1.285 0.870 1.515 ;
        RECT  0.850 1.930 1.490 2.050 ;
        RECT  1.490 1.425 1.610 2.050 ;
        RECT  1.610 1.425 1.700 1.550 ;
        RECT  1.700 1.040 1.860 1.550 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.255 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.160 0.300 ;
        RECT  1.160 -0.300 1.380 0.340 ;
        RECT  1.380 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.140 1.410 1.240 1.810 ;
        RECT  1.140 0.470 2.260 0.590 ;
        RECT  2.260 0.470 2.380 1.000 ;
        RECT  2.380 0.880 2.660 1.000 ;
        RECT  2.660 0.880 2.820 1.150 ;
        RECT  1.780 0.710 2.020 0.870 ;
        RECT  2.020 0.710 2.140 2.020 ;
        RECT  2.140 1.170 2.510 1.330 ;
        RECT  0.210 1.470 0.250 1.710 ;
        RECT  0.210 0.420 0.250 0.960 ;
        RECT  0.250 0.800 0.790 0.960 ;
        RECT  1.020 0.470 1.140 1.810 ;
        RECT  0.995 0.470 1.020 0.590 ;
        RECT  0.750 0.430 0.995 0.590 ;
        RECT  1.730 1.860 2.020 2.020 ;
        RECT  0.090 0.420 0.210 1.710 ;
    END
END BUFTD2

MACRO BUFTD20
    CLASS CORE ;
    FOREIGN BUFTD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  5.290 1.860 6.000 2.020 ;
        RECT  6.000 1.640 8.270 2.020 ;
        RECT  5.100 0.480 8.270 0.640 ;
        RECT  8.270 0.480 8.690 2.020 ;
        RECT  8.690 1.640 11.740 2.020 ;
        RECT  8.690 0.480 11.760 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.040 0.410 1.260 ;
        RECT  0.410 0.470 0.530 1.260 ;
        RECT  0.530 0.470 2.650 0.590 ;
        RECT  2.650 0.470 2.790 0.845 ;
        RECT  2.790 0.725 3.290 0.845 ;
        RECT  3.290 0.725 3.410 1.235 ;
        RECT  3.410 1.005 3.750 1.235 ;
        RECT  3.410 0.725 4.480 0.845 ;
        RECT  4.480 0.725 4.640 1.220 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.095 2.330 1.255 ;
        RECT  2.330 1.005 2.710 1.255 ;
        RECT  2.710 1.005 2.790 1.480 ;
        RECT  2.790 1.095 2.870 1.480 ;
        RECT  2.870 1.360 3.880 1.480 ;
        RECT  3.880 1.080 4.040 1.480 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.710 0.300 ;
        RECT  4.710 -0.300 4.930 0.340 ;
        RECT  4.930 -0.300 5.510 0.300 ;
        RECT  5.510 -0.300 5.730 0.340 ;
        RECT  5.730 -0.300 6.300 0.300 ;
        RECT  6.300 -0.300 6.520 0.340 ;
        RECT  6.520 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.650 1.020 0.790 1.510 ;
        RECT  0.250 1.390 0.650 1.510 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.210 0.420 0.250 0.900 ;
        RECT  0.210 1.390 0.250 2.100 ;
        RECT  0.090 0.420 0.210 2.100 ;
        RECT  4.890 1.170 5.420 1.330 ;
        RECT  4.880 1.170 4.890 1.810 ;
        RECT  4.760 0.470 4.880 1.810 ;
        RECT  4.570 0.470 4.760 0.590 ;
        RECT  2.580 1.650 4.760 1.810 ;
        RECT  4.350 0.430 4.570 0.590 ;
        RECT  3.380 0.470 4.350 0.590 ;
        RECT  5.570 0.890 5.730 1.620 ;
        RECT  5.130 1.500 5.570 1.620 ;
        RECT  5.010 1.500 5.130 2.050 ;
        RECT  2.450 1.930 5.010 2.050 ;
        RECT  2.290 1.430 2.450 2.050 ;
        RECT  1.040 0.710 2.420 0.870 ;
        RECT  1.260 1.430 2.290 1.550 ;
        RECT  1.100 1.430 1.260 1.930 ;
        RECT  1.040 1.430 1.100 1.550 ;
        RECT  0.920 0.710 1.040 1.550 ;
        RECT  0.760 0.710 0.920 0.870 ;
        RECT  3.140 0.430 3.380 0.590 ;
        RECT  0.060 1.960 0.090 2.100 ;
        LAYER M1 ;
        RECT  6.000 1.640 8.055 2.020 ;
        RECT  5.100 0.480 8.055 0.640 ;
        RECT  5.290 1.860 6.000 2.020 ;
        RECT  8.905 0.480 11.760 0.640 ;
        RECT  8.905 1.640 11.740 2.020 ;
    END
END BUFTD20

MACRO BUFTD24
    CLASS CORE ;
    FOREIGN BUFTD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  5.300 1.860 6.010 2.020 ;
        RECT  6.010 1.640 8.270 2.020 ;
        RECT  5.110 0.480 8.270 0.640 ;
        RECT  8.270 0.480 8.690 2.020 ;
        RECT  8.690 1.640 13.320 2.020 ;
        RECT  8.690 0.480 13.340 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.040 0.410 1.260 ;
        RECT  0.410 0.470 0.530 1.260 ;
        RECT  0.530 0.470 2.650 0.590 ;
        RECT  2.650 0.470 2.790 0.845 ;
        RECT  2.790 0.725 3.290 0.845 ;
        RECT  3.290 0.725 3.410 1.235 ;
        RECT  3.410 1.005 3.750 1.235 ;
        RECT  3.410 0.725 4.480 0.845 ;
        RECT  4.480 0.725 4.640 1.220 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.095 2.330 1.255 ;
        RECT  2.330 1.005 2.710 1.255 ;
        RECT  2.710 1.005 2.790 1.480 ;
        RECT  2.790 1.095 2.870 1.480 ;
        RECT  2.870 1.360 3.880 1.480 ;
        RECT  3.880 1.080 4.040 1.480 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.940 0.340 ;
        RECT  4.940 -0.300 5.520 0.300 ;
        RECT  5.520 -0.300 5.740 0.340 ;
        RECT  5.740 -0.300 6.310 0.300 ;
        RECT  6.310 -0.300 6.530 0.340 ;
        RECT  6.530 -0.300 13.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 13.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.650 1.020 0.790 1.510 ;
        RECT  0.250 1.390 0.650 1.510 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.210 0.420 0.250 0.900 ;
        RECT  0.210 1.390 0.250 2.100 ;
        RECT  0.090 0.420 0.210 2.100 ;
        RECT  4.890 1.170 5.430 1.330 ;
        RECT  4.880 1.170 4.890 1.810 ;
        RECT  4.760 0.470 4.880 1.810 ;
        RECT  4.570 0.470 4.760 0.590 ;
        RECT  2.580 1.650 4.760 1.810 ;
        RECT  4.350 0.430 4.570 0.590 ;
        RECT  3.380 0.470 4.350 0.590 ;
        RECT  5.580 0.890 5.740 1.620 ;
        RECT  5.130 1.500 5.580 1.620 ;
        RECT  5.010 1.500 5.130 2.050 ;
        RECT  2.450 1.930 5.010 2.050 ;
        RECT  2.290 1.430 2.450 2.050 ;
        RECT  1.040 0.710 2.420 0.870 ;
        RECT  1.260 1.430 2.290 1.550 ;
        RECT  1.100 1.430 1.260 1.930 ;
        RECT  1.040 1.430 1.100 1.550 ;
        RECT  0.920 0.710 1.040 1.550 ;
        RECT  3.140 0.430 3.380 0.590 ;
        RECT  0.060 1.960 0.090 2.100 ;
        RECT  0.760 0.710 0.920 0.870 ;
        LAYER M1 ;
        RECT  6.010 1.640 8.055 2.020 ;
        RECT  5.110 0.480 8.055 0.640 ;
        RECT  5.300 1.860 6.010 2.020 ;
        RECT  8.905 0.480 13.340 0.640 ;
        RECT  8.905 1.640 13.320 2.020 ;
    END
END BUFTD24

MACRO BUFTD3
    CLASS CORE ;
    FOREIGN BUFTD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.510 1.640 2.830 2.020 ;
        RECT  2.830 1.425 3.130 2.020 ;
        RECT  2.510 0.500 3.130 0.660 ;
        RECT  3.130 0.500 3.250 2.020 ;
        RECT  3.250 1.640 3.460 2.020 ;
        RECT  3.250 0.500 3.460 0.660 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.110 0.410 1.330 ;
        RECT  0.410 1.110 0.550 1.515 ;
        RECT  0.550 1.285 0.710 1.515 ;
        RECT  0.710 1.285 0.850 2.050 ;
        RECT  0.850 1.285 0.870 1.515 ;
        RECT  0.850 1.930 1.550 2.050 ;
        RECT  1.550 1.425 1.670 2.050 ;
        RECT  1.670 1.425 1.750 1.550 ;
        RECT  1.750 1.000 1.910 1.550 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.255 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 1.380 2.820 ;
        RECT  1.380 2.180 1.600 2.820 ;
        RECT  1.600 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.020 0.470 1.140 1.810 ;
        RECT  1.140 1.410 1.240 1.810 ;
        RECT  1.140 0.470 2.270 0.590 ;
        RECT  2.270 0.470 2.390 1.000 ;
        RECT  2.390 0.880 2.670 1.000 ;
        RECT  2.670 0.880 2.830 1.150 ;
        RECT  1.830 0.710 2.030 0.870 ;
        RECT  2.030 0.710 2.150 2.020 ;
        RECT  2.150 1.170 2.520 1.330 ;
        RECT  0.210 1.470 0.250 1.710 ;
        RECT  0.210 0.420 0.250 0.960 ;
        RECT  0.250 0.800 0.790 0.960 ;
        RECT  0.995 0.470 1.020 0.590 ;
        RECT  1.790 1.860 2.030 2.020 ;
        RECT  0.090 0.420 0.210 1.710 ;
        RECT  0.750 0.430 0.995 0.590 ;
        LAYER M1 ;
        RECT  2.510 0.500 3.130 0.660 ;
        RECT  2.510 1.640 2.615 2.020 ;
        RECT  3.130 0.500 3.250 1.255 ;
        RECT  3.250 0.500 3.460 0.660 ;
    END
END BUFTD3

MACRO BUFTD4
    CLASS CORE ;
    FOREIGN BUFTD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.640 3.150 2.020 ;
        RECT  2.500 0.500 3.150 0.660 ;
        RECT  3.150 0.500 3.570 2.020 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.110 0.410 1.330 ;
        RECT  0.410 1.110 0.550 1.515 ;
        RECT  0.550 1.285 0.710 1.515 ;
        RECT  0.710 1.285 0.850 2.050 ;
        RECT  0.850 1.285 0.870 1.515 ;
        RECT  0.850 1.930 1.550 2.050 ;
        RECT  1.550 1.425 1.670 2.050 ;
        RECT  1.670 1.425 1.740 1.550 ;
        RECT  1.740 0.980 1.900 1.550 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.255 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 1.380 2.820 ;
        RECT  1.380 2.180 1.600 2.820 ;
        RECT  1.600 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.020 0.710 2.140 1.830 ;
        RECT  2.140 1.170 2.520 1.330 ;
        RECT  0.210 1.470 0.250 1.710 ;
        RECT  0.210 0.420 0.250 0.960 ;
        RECT  0.250 0.800 0.790 0.960 ;
        RECT  1.840 0.710 2.020 0.860 ;
        RECT  2.010 1.670 2.020 1.830 ;
        RECT  2.670 0.880 2.830 1.150 ;
        RECT  2.380 0.880 2.670 1.000 ;
        RECT  2.260 0.470 2.380 1.000 ;
        RECT  1.140 0.470 2.260 0.590 ;
        RECT  1.140 1.410 1.240 1.810 ;
        RECT  1.020 0.470 1.140 1.810 ;
        RECT  0.995 0.470 1.020 0.590 ;
        RECT  0.750 0.430 0.995 0.590 ;
        RECT  1.790 1.670 2.010 2.090 ;
        RECT  0.090 0.420 0.210 1.710 ;
        LAYER M1 ;
        RECT  2.500 0.500 2.935 0.660 ;
        RECT  2.490 1.640 2.935 2.020 ;
    END
END BUFTD4

MACRO BUFTD6
    CLASS CORE ;
    FOREIGN BUFTD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.390 1.640 4.110 2.020 ;
        RECT  3.390 0.480 4.110 0.640 ;
        RECT  4.110 0.480 4.530 2.020 ;
        RECT  4.530 1.640 5.020 2.020 ;
        RECT  4.530 0.480 5.040 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.030 0.490 2.050 ;
        RECT  0.490 1.930 1.700 2.050 ;
        RECT  1.700 1.395 1.820 2.050 ;
        RECT  1.820 1.395 2.330 1.515 ;
        RECT  2.330 1.005 2.450 1.515 ;
        RECT  2.450 1.005 2.790 1.235 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.880 1.510 1.810 ;
        RECT  1.105 0.880 1.390 1.040 ;
        RECT  0.745 1.690 1.390 1.810 ;
        RECT  0.625 0.790 0.745 1.810 ;
        RECT  0.250 0.790 0.625 0.910 ;
        RECT  0.230 0.420 0.250 0.910 ;
        RECT  3.270 0.940 3.500 1.090 ;
        RECT  3.150 0.470 3.270 1.090 ;
        RECT  1.680 0.470 3.150 0.590 ;
        RECT  1.460 0.430 1.680 0.590 ;
        RECT  0.990 0.470 1.460 0.590 ;
        RECT  0.985 1.410 1.260 1.570 ;
        RECT  0.985 0.430 0.990 0.590 ;
        RECT  0.865 0.430 0.985 1.570 ;
        RECT  3.620 1.170 3.860 1.330 ;
        RECT  3.030 1.210 3.620 1.330 ;
        RECT  2.910 0.710 3.030 1.770 ;
        RECT  2.890 1.960 2.920 2.100 ;
        RECT  2.395 0.710 2.910 0.870 ;
        RECT  2.890 1.650 2.910 1.770 ;
        RECT  2.730 1.650 2.890 2.100 ;
        RECT  2.700 1.930 2.730 2.100 ;
        RECT  2.220 1.930 2.700 2.050 ;
        RECT  2.190 1.930 2.220 2.090 ;
        RECT  2.030 1.640 2.190 2.090 ;
        RECT  2.000 1.930 2.030 2.090 ;
        RECT  0.750 0.430 0.865 0.590 ;
        RECT  0.090 0.420 0.230 1.710 ;
        LAYER M1 ;
        RECT  4.745 1.640 5.020 2.020 ;
        RECT  4.745 0.480 5.040 0.640 ;
        RECT  3.390 1.640 3.895 2.020 ;
        RECT  3.390 0.480 3.895 0.640 ;
    END
END BUFTD6

MACRO BUFTD8
    CLASS CORE ;
    FOREIGN BUFTD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.640 4.430 2.020 ;
        RECT  3.350 0.480 4.430 0.640 ;
        RECT  4.430 0.480 4.850 2.020 ;
        RECT  4.850 1.640 5.660 2.020 ;
        RECT  4.850 0.480 5.680 0.640 ;
        END
    END Z
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.030 0.490 2.050 ;
        RECT  0.490 1.930 1.700 2.050 ;
        RECT  1.700 1.395 1.820 2.050 ;
        RECT  1.820 1.395 2.320 1.515 ;
        RECT  2.320 1.005 2.480 1.515 ;
        END
    END OE
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.880 1.510 1.810 ;
        RECT  1.105 0.880 1.390 1.040 ;
        RECT  0.745 1.690 1.390 1.810 ;
        RECT  0.625 0.790 0.745 1.810 ;
        RECT  0.250 0.790 0.625 0.910 ;
        RECT  0.230 0.430 0.250 0.910 ;
        RECT  3.180 0.940 3.480 1.090 ;
        RECT  3.060 0.470 3.180 1.090 ;
        RECT  1.680 0.470 3.060 0.590 ;
        RECT  1.460 0.430 1.680 0.590 ;
        RECT  0.990 0.470 1.460 0.590 ;
        RECT  0.985 1.410 1.260 1.570 ;
        RECT  0.985 0.430 0.990 0.590 ;
        RECT  0.865 0.430 0.985 1.570 ;
        RECT  3.600 1.170 3.840 1.330 ;
        RECT  2.870 1.210 3.600 1.330 ;
        RECT  2.870 1.960 2.900 2.100 ;
        RECT  2.710 0.710 2.870 2.100 ;
        RECT  2.405 0.710 2.710 0.870 ;
        RECT  2.680 1.930 2.710 2.100 ;
        RECT  2.210 1.930 2.680 2.050 ;
        RECT  2.180 1.930 2.210 2.090 ;
        RECT  2.020 1.640 2.180 2.090 ;
        RECT  1.990 1.930 2.020 2.090 ;
        RECT  0.750 0.430 0.865 0.590 ;
        RECT  0.090 0.430 0.230 1.690 ;
        LAYER M1 ;
        RECT  3.350 0.480 4.215 0.640 ;
        RECT  3.370 1.640 4.215 2.020 ;
        RECT  5.065 0.480 5.680 0.640 ;
        RECT  5.065 1.640 5.660 2.020 ;
    END
END BUFTD8

MACRO CKAN2D0
    CLASS CORE ;
    FOREIGN CKAN2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 0.620 1.350 0.840 ;
        RECT  1.350 0.620 1.510 1.890 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.850 0.300 ;
        RECT  0.850 -0.300 1.070 0.340 ;
        RECT  1.070 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.920 2.820 ;
        RECT  0.920 2.180 1.140 2.820 ;
        RECT  1.140 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.010 0.650 1.170 1.660 ;
        RECT  0.160 0.650 1.010 0.810 ;
        RECT  0.490 1.500 1.010 1.660 ;
    END
END CKAN2D0

MACRO CKAN2D1
    CLASS CORE ;
    FOREIGN CKAN2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.350 0.600 1.510 2.100 ;
        RECT  1.510 1.960 1.540 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.100 0.340 ;
        RECT  1.100 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.920 2.820 ;
        RECT  0.920 2.180 1.140 2.820 ;
        RECT  1.140 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.650 1.230 1.660 ;
        RECT  0.160 0.650 1.070 0.810 ;
        RECT  0.490 1.500 1.070 1.660 ;
    END
END CKAN2D1

MACRO CKAN2D2
    CLASS CORE ;
    FOREIGN CKAN2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.960 1.280 2.100 ;
        RECT  1.280 1.390 1.370 2.100 ;
        RECT  1.280 0.420 1.370 0.920 ;
        RECT  1.370 0.420 1.440 2.100 ;
        RECT  1.440 1.960 1.470 2.100 ;
        RECT  1.440 0.800 1.510 1.515 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.840 0.300 ;
        RECT  0.840 -0.300 1.060 0.340 ;
        RECT  1.060 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.860 2.820 ;
        RECT  0.860 2.180 1.080 2.820 ;
        RECT  1.080 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.690 1.160 1.510 ;
        RECT  0.150 0.690 1.000 0.850 ;
        RECT  0.660 1.390 1.000 1.510 ;
        RECT  0.500 1.390 0.660 1.890 ;
    END
END CKAN2D2

MACRO CKAN2D4
    CLASS CORE ;
    FOREIGN CKAN2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.640 1.870 2.020 ;
        RECT  1.240 0.500 1.870 0.880 ;
        RECT  1.870 0.500 2.290 2.020 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.240 ;
        RECT  0.550 1.080 0.770 1.240 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.790 0.300 ;
        RECT  0.790 -0.300 1.010 0.340 ;
        RECT  1.010 -0.300 1.660 0.300 ;
        RECT  1.660 -0.300 1.880 0.340 ;
        RECT  1.880 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.020 1.080 1.580 1.240 ;
        RECT  0.900 0.470 1.020 1.510 ;
        RECT  0.290 0.470 0.900 0.590 ;
        RECT  0.620 1.390 0.900 1.510 ;
        RECT  0.460 1.390 0.620 1.890 ;
        RECT  0.070 0.470 0.290 0.885 ;
        LAYER M1 ;
        RECT  1.140 1.640 1.655 2.020 ;
        RECT  1.240 0.500 1.655 0.880 ;
    END
END CKAN2D4

MACRO CKAN2D8
    CLASS CORE ;
    FOREIGN CKAN2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.640 2.830 2.020 ;
        RECT  1.880 0.500 2.830 0.880 ;
        RECT  2.830 0.500 3.250 2.020 ;
        RECT  3.250 1.640 4.270 2.020 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.320 1.515 ;
        RECT  1.320 1.030 1.480 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.470 0.300 ;
        RECT  1.470 -0.300 1.690 0.340 ;
        RECT  1.690 -0.300 2.300 0.300 ;
        RECT  2.300 -0.300 2.520 0.340 ;
        RECT  2.520 -0.300 3.120 0.300 ;
        RECT  3.120 -0.300 3.340 0.340 ;
        RECT  3.340 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.450 2.820 ;
        RECT  4.450 2.180 4.670 2.820 ;
        RECT  4.670 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.740 1.080 2.490 1.240 ;
        RECT  1.620 0.725 1.740 1.790 ;
        RECT  0.780 0.725 1.620 0.885 ;
        RECT  0.420 1.635 1.620 1.790 ;
        LAYER M1 ;
        RECT  1.860 1.640 2.615 2.020 ;
        RECT  1.880 0.500 2.615 0.880 ;
        RECT  3.465 1.640 4.270 2.020 ;
    END
END CKAN2D8

MACRO CKBD0
    CLASS CORE ;
    FOREIGN CKBD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.985 0.240 1.515 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.430 1.190 1.925 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.340 ;
        RECT  0.760 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 2.180 0.760 2.820 ;
        RECT  0.760 2.220 1.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.480 0.910 1.795 ;
        RECT  0.100 1.635 0.750 1.795 ;
        RECT  0.100 0.480 0.750 0.640 ;
    END
END CKBD0

MACRO CKBD1
    CLASS CORE ;
    FOREIGN CKBD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.350 0.420 1.510 2.100 ;
        RECT  1.510 1.960 1.540 2.100 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.860 0.300 ;
        RECT  0.860 -0.300 1.080 0.340 ;
        RECT  1.080 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.860 2.820 ;
        RECT  0.860 2.180 1.080 2.820 ;
        RECT  1.080 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.630 1.080 1.230 1.240 ;
        RECT  0.630 1.960 0.660 2.100 ;
        RECT  0.470 0.420 0.630 2.100 ;
        RECT  0.440 1.960 0.470 2.100 ;
    END
END CKBD1

MACRO CKBD12
    CLASS CORE ;
    FOREIGN CKBD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.440 1.650 4.110 2.030 ;
        RECT  2.890 0.470 4.110 0.710 ;
        RECT  4.110 0.470 4.530 2.030 ;
        RECT  4.530 1.650 6.320 2.030 ;
        RECT  4.530 0.470 6.330 0.710 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.510 0.300 ;
        RECT  2.510 -0.300 2.730 0.340 ;
        RECT  2.730 -0.300 3.310 0.300 ;
        RECT  3.310 -0.300 3.530 0.340 ;
        RECT  3.530 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.340 ;
        RECT  4.330 -0.300 4.910 0.300 ;
        RECT  4.910 -0.300 5.130 0.340 ;
        RECT  5.130 -0.300 5.710 0.300 ;
        RECT  5.710 -0.300 5.930 0.340 ;
        RECT  5.930 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.680 2.820 ;
        RECT  5.680 2.180 5.900 2.820 ;
        RECT  5.900 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.880 3.860 1.040 ;
        RECT  2.190 0.450 2.350 1.040 ;
        RECT  1.990 0.885 2.190 1.040 ;
        RECT  1.990 1.960 2.020 2.100 ;
        RECT  1.830 0.885 1.990 2.100 ;
        RECT  1.630 0.885 1.830 1.045 ;
        RECT  1.800 1.960 1.830 2.100 ;
        RECT  1.470 0.450 1.630 1.045 ;
        RECT  1.300 0.885 1.470 1.045 ;
        RECT  1.300 1.960 1.330 2.100 ;
        RECT  1.140 0.885 1.300 2.100 ;
        RECT  0.910 0.885 1.140 1.045 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  0.750 0.450 0.910 1.045 ;
        RECT  0.610 0.885 0.750 1.045 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 0.885 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  2.890 0.470 3.895 0.710 ;
        RECT  4.745 0.470 6.330 0.710 ;
        RECT  4.745 1.650 6.320 2.030 ;
        RECT  2.440 1.650 3.895 2.030 ;
    END
END CKBD12

MACRO CKBD16
    CLASS CORE ;
    FOREIGN CKBD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.650 5.070 2.030 ;
        RECT  3.230 0.470 5.070 0.710 ;
        RECT  5.070 0.470 5.490 2.030 ;
        RECT  5.490 0.470 7.490 0.710 ;
        RECT  5.490 1.650 7.880 2.030 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.420 0.300 ;
        RECT  0.420 -0.300 0.640 0.340 ;
        RECT  0.640 -0.300 1.240 0.300 ;
        RECT  1.240 -0.300 1.460 0.340 ;
        RECT  1.460 -0.300 2.050 0.300 ;
        RECT  2.050 -0.300 2.270 0.340 ;
        RECT  2.270 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.650 0.300 ;
        RECT  3.650 -0.300 3.870 0.340 ;
        RECT  3.870 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 5.250 0.300 ;
        RECT  5.250 -0.300 5.470 0.340 ;
        RECT  5.470 -0.300 6.050 0.300 ;
        RECT  6.050 -0.300 6.270 0.340 ;
        RECT  6.270 -0.300 6.850 0.300 ;
        RECT  6.850 -0.300 7.070 0.340 ;
        RECT  7.070 -0.300 7.650 0.300 ;
        RECT  7.650 -0.300 7.870 0.340 ;
        RECT  7.870 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.240 2.820 ;
        RECT  7.240 2.180 7.460 2.820 ;
        RECT  7.460 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.730 0.880 4.745 1.040 ;
        RECT  2.730 1.960 2.760 2.100 ;
        RECT  2.640 0.880 2.730 2.100 ;
        RECT  2.570 0.420 2.640 2.100 ;
        RECT  2.480 0.420 2.570 1.040 ;
        RECT  2.540 1.960 2.570 2.100 ;
        RECT  2.020 0.880 2.480 1.040 ;
        RECT  2.020 1.960 2.050 2.100 ;
        RECT  1.860 0.880 2.020 2.100 ;
        RECT  1.840 0.880 1.860 1.040 ;
        RECT  1.830 1.960 1.860 2.100 ;
        RECT  1.680 0.420 1.840 1.040 ;
        RECT  1.320 0.880 1.680 1.040 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.160 0.880 1.320 2.100 ;
        RECT  1.020 0.880 1.160 1.040 ;
        RECT  1.130 1.960 1.160 2.100 ;
        RECT  0.860 0.420 1.020 1.040 ;
        RECT  0.620 0.880 0.860 1.040 ;
        RECT  0.620 1.960 0.650 2.100 ;
        RECT  0.460 0.880 0.620 2.100 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  3.230 0.470 4.855 0.710 ;
        RECT  5.705 0.470 7.490 0.710 ;
        RECT  5.705 1.650 7.880 2.030 ;
        RECT  3.180 1.650 4.855 2.030 ;
    END
END CKBD16

MACRO CKBD2
    CLASS CORE ;
    FOREIGN CKBD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.960 0.890 2.100 ;
        RECT  0.890 1.390 1.050 2.100 ;
        RECT  1.050 1.960 1.080 2.100 ;
        RECT  1.050 1.390 1.350 1.515 ;
        RECT  1.350 0.420 1.510 1.515 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.870 0.300 ;
        RECT  0.870 -0.300 1.090 0.340 ;
        RECT  1.090 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.100 1.390 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.260 1.390 0.480 1.510 ;
        RECT  0.480 0.460 0.600 1.510 ;
        RECT  0.600 0.460 0.640 1.240 ;
        RECT  0.640 1.080 1.230 1.240 ;
        RECT  0.070 1.960 0.100 2.100 ;
    END
END CKBD2

MACRO CKBD20
    CLASS CORE ;
    FOREIGN CKBD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.020 1.650 6.670 2.030 ;
        RECT  3.890 0.470 6.670 0.695 ;
        RECT  6.670 0.470 7.090 2.030 ;
        RECT  7.090 1.650 9.700 2.030 ;
        RECT  7.090 0.470 9.730 0.695 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.400 0.300 ;
        RECT  0.400 -0.300 0.620 0.340 ;
        RECT  0.620 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 1.960 0.300 ;
        RECT  1.960 -0.300 2.180 0.340 ;
        RECT  2.180 -0.300 2.740 0.300 ;
        RECT  2.740 -0.300 2.960 0.340 ;
        RECT  2.960 -0.300 3.520 0.300 ;
        RECT  3.520 -0.300 3.740 0.340 ;
        RECT  3.740 -0.300 4.300 0.300 ;
        RECT  4.300 -0.300 4.520 0.340 ;
        RECT  4.520 -0.300 5.090 0.300 ;
        RECT  5.090 -0.300 5.310 0.340 ;
        RECT  5.310 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.340 ;
        RECT  6.110 -0.300 6.690 0.300 ;
        RECT  6.690 -0.300 6.910 0.340 ;
        RECT  6.910 -0.300 7.490 0.300 ;
        RECT  7.490 -0.300 7.710 0.340 ;
        RECT  7.710 -0.300 8.290 0.300 ;
        RECT  8.290 -0.300 8.510 0.340 ;
        RECT  8.510 -0.300 9.090 0.300 ;
        RECT  9.090 -0.300 9.310 0.340 ;
        RECT  9.310 -0.300 9.890 0.300 ;
        RECT  9.890 -0.300 10.110 0.340 ;
        RECT  10.110 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.630 2.820 ;
        RECT  3.630 2.180 3.850 2.820 ;
        RECT  3.850 2.220 4.410 2.820 ;
        RECT  4.410 2.180 4.630 2.820 ;
        RECT  4.630 2.220 5.190 2.820 ;
        RECT  5.190 2.180 5.410 2.820 ;
        RECT  5.410 2.220 5.970 2.820 ;
        RECT  5.970 2.180 6.190 2.820 ;
        RECT  6.190 2.220 6.750 2.820 ;
        RECT  6.750 2.180 6.970 2.820 ;
        RECT  6.970 2.220 7.530 2.820 ;
        RECT  7.530 2.180 7.750 2.820 ;
        RECT  7.750 2.220 8.310 2.820 ;
        RECT  8.310 2.180 8.530 2.820 ;
        RECT  8.530 2.220 9.090 2.820 ;
        RECT  9.090 2.180 9.310 2.820 ;
        RECT  9.310 2.220 9.880 2.820 ;
        RECT  9.880 2.180 10.100 2.820 ;
        RECT  10.100 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.420 0.865 5.055 1.025 ;
        RECT  3.420 1.960 3.450 2.100 ;
        RECT  3.320 0.865 3.420 2.100 ;
        RECT  3.260 0.420 3.320 2.100 ;
        RECT  3.160 0.420 3.260 1.005 ;
        RECT  3.230 1.960 3.260 2.100 ;
        RECT  2.720 0.845 3.160 1.005 ;
        RECT  2.720 1.960 2.750 2.100 ;
        RECT  2.560 0.845 2.720 2.100 ;
        RECT  2.540 0.845 2.560 1.005 ;
        RECT  2.530 1.960 2.560 2.100 ;
        RECT  2.380 0.420 2.540 1.005 ;
        RECT  2.020 0.845 2.380 1.005 ;
        RECT  2.020 1.960 2.050 2.100 ;
        RECT  1.860 0.845 2.020 2.100 ;
        RECT  1.760 0.845 1.860 1.005 ;
        RECT  1.830 1.960 1.860 2.100 ;
        RECT  1.600 0.420 1.760 1.005 ;
        RECT  1.320 0.845 1.600 1.005 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.160 0.845 1.320 2.100 ;
        RECT  0.980 0.845 1.160 1.005 ;
        RECT  1.130 1.960 1.160 2.100 ;
        RECT  0.820 0.420 0.980 1.005 ;
        RECT  0.620 0.845 0.820 1.005 ;
        RECT  0.620 1.960 0.650 2.100 ;
        RECT  0.460 0.845 0.620 2.100 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  3.890 0.470 6.455 0.695 ;
        RECT  7.755 0.470 9.730 0.695 ;
        RECT  7.305 1.650 9.700 2.030 ;
        RECT  4.020 1.650 6.455 2.030 ;
    END
END CKBD20

MACRO CKBD24
    CLASS CORE ;
    FOREIGN CKBD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.690 1.650 7.630 2.030 ;
        RECT  4.530 0.470 7.630 0.710 ;
        RECT  7.630 0.470 8.050 2.030 ;
        RECT  8.050 1.650 10.520 2.030 ;
        RECT  8.050 0.470 11.030 0.710 ;
        RECT  10.520 1.650 11.320 1.810 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.830 0.300 ;
        RECT  0.830 -0.300 1.050 0.340 ;
        RECT  1.050 -0.300 1.660 0.300 ;
        RECT  1.660 -0.300 1.880 0.340 ;
        RECT  1.880 -0.300 2.490 0.300 ;
        RECT  2.490 -0.300 2.710 0.340 ;
        RECT  2.710 -0.300 3.320 0.300 ;
        RECT  3.320 -0.300 3.540 0.340 ;
        RECT  3.540 -0.300 4.140 0.300 ;
        RECT  4.140 -0.300 4.360 0.340 ;
        RECT  4.360 -0.300 4.940 0.300 ;
        RECT  4.940 -0.300 5.160 0.340 ;
        RECT  5.160 -0.300 5.720 0.300 ;
        RECT  5.720 -0.300 5.940 0.340 ;
        RECT  5.940 -0.300 6.500 0.300 ;
        RECT  6.500 -0.300 6.720 0.340 ;
        RECT  6.720 -0.300 7.280 0.300 ;
        RECT  7.280 -0.300 7.500 0.340 ;
        RECT  7.500 -0.300 8.060 0.300 ;
        RECT  8.060 -0.300 8.280 0.340 ;
        RECT  8.280 -0.300 8.840 0.300 ;
        RECT  8.840 -0.300 9.060 0.340 ;
        RECT  9.060 -0.300 9.620 0.300 ;
        RECT  9.620 -0.300 9.840 0.340 ;
        RECT  9.840 -0.300 10.400 0.300 ;
        RECT  10.400 -0.300 10.620 0.340 ;
        RECT  10.620 -0.300 11.180 0.300 ;
        RECT  11.180 -0.300 11.400 0.340 ;
        RECT  11.400 -0.300 11.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 10.690 2.820 ;
        RECT  10.690 2.180 10.910 2.820 ;
        RECT  10.910 2.220 11.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.120 0.880 5.730 1.040 ;
        RECT  4.120 1.960 4.150 2.100 ;
        RECT  3.960 0.880 4.120 2.100 ;
        RECT  3.920 0.880 3.960 1.040 ;
        RECT  3.930 1.960 3.960 2.100 ;
        RECT  3.760 0.420 3.920 1.040 ;
        RECT  3.420 0.880 3.760 1.040 ;
        RECT  3.420 1.960 3.450 2.100 ;
        RECT  3.260 0.880 3.420 2.100 ;
        RECT  3.090 0.880 3.260 1.040 ;
        RECT  3.230 1.960 3.260 2.100 ;
        RECT  2.930 0.420 3.090 1.040 ;
        RECT  2.720 0.880 2.930 1.040 ;
        RECT  2.720 1.960 2.750 2.100 ;
        RECT  2.560 0.880 2.720 2.100 ;
        RECT  2.260 0.880 2.560 1.040 ;
        RECT  2.530 1.960 2.560 2.100 ;
        RECT  2.100 0.420 2.260 1.040 ;
        RECT  2.020 0.880 2.100 1.040 ;
        RECT  2.020 1.960 2.050 2.100 ;
        RECT  1.860 0.880 2.020 2.100 ;
        RECT  1.430 0.880 1.860 1.040 ;
        RECT  1.830 1.960 1.860 2.100 ;
        RECT  1.320 0.420 1.430 1.040 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.270 0.420 1.320 2.100 ;
        RECT  1.160 0.880 1.270 2.100 ;
        RECT  0.620 0.880 1.160 1.040 ;
        RECT  1.130 1.960 1.160 2.100 ;
        RECT  0.620 1.960 0.650 2.100 ;
        RECT  0.600 0.880 0.620 2.100 ;
        RECT  0.460 0.420 0.600 2.100 ;
        RECT  0.440 0.420 0.460 1.040 ;
        RECT  0.430 1.960 0.460 2.100 ;
        LAYER M1 ;
        RECT  10.520 1.650 11.320 1.810 ;
        RECT  8.265 0.470 11.030 0.710 ;
        RECT  4.530 0.470 7.415 0.710 ;
        RECT  8.265 1.650 10.520 2.030 ;
        RECT  4.690 1.650 7.415 2.030 ;
    END
END CKBD24

MACRO CKBD3
    CLASS CORE ;
    FOREIGN CKBD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.640 1.550 2.020 ;
        RECT  1.550 0.500 1.970 2.020 ;
        RECT  1.970 1.640 2.180 2.020 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.960 1.080 1.320 1.240 ;
        RECT  0.800 0.420 0.960 1.240 ;
        RECT  0.660 1.080 0.800 1.240 ;
        RECT  0.660 1.960 0.690 2.100 ;
        RECT  0.500 1.080 0.660 2.100 ;
        RECT  0.470 1.960 0.500 2.100 ;
        LAYER M1 ;
        RECT  1.210 1.640 1.335 2.020 ;
    END
END CKBD3

MACRO CKBD4
    CLASS CORE ;
    FOREIGN CKBD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.640 1.550 2.020 ;
        RECT  1.520 0.480 1.550 0.620 ;
        RECT  1.550 0.480 1.970 2.020 ;
        RECT  1.970 1.640 2.120 2.020 ;
        RECT  1.970 0.480 2.500 0.640 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 1.070 1.270 1.230 ;
        RECT  0.790 0.420 0.950 1.230 ;
        RECT  0.630 1.070 0.790 1.230 ;
        RECT  0.630 1.960 0.660 2.100 ;
        RECT  0.470 1.070 0.630 2.100 ;
        RECT  0.440 1.960 0.470 2.100 ;
        LAYER M1 ;
        RECT  1.160 1.640 1.335 2.020 ;
        RECT  2.185 0.480 2.500 0.640 ;
    END
END CKBD4

MACRO CKBD6
    CLASS CORE ;
    FOREIGN CKBD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.255 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.470 1.640 2.190 2.020 ;
        RECT  1.600 0.550 2.190 0.710 ;
        RECT  2.190 0.550 2.610 2.020 ;
        RECT  2.610 1.640 3.090 2.020 ;
        RECT  2.610 0.550 3.460 0.710 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.410 0.300 ;
        RECT  0.410 -0.300 0.630 0.340 ;
        RECT  0.630 -0.300 1.220 0.300 ;
        RECT  1.220 -0.300 1.440 0.340 ;
        RECT  1.440 -0.300 2.030 0.300 ;
        RECT  2.030 -0.300 2.250 0.340 ;
        RECT  2.250 -0.300 2.830 0.300 ;
        RECT  2.830 -0.300 3.050 0.340 ;
        RECT  3.050 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 1.045 1.840 1.205 ;
        RECT  0.950 0.460 1.000 1.205 ;
        RECT  0.950 1.960 0.980 2.100 ;
        RECT  0.840 0.460 0.950 2.100 ;
        RECT  0.790 1.045 0.840 2.100 ;
        RECT  0.250 1.390 0.790 1.510 ;
        RECT  0.760 1.960 0.790 2.100 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.090 1.390 0.250 2.100 ;
        RECT  0.060 1.960 0.090 2.100 ;
        LAYER M1 ;
        RECT  1.470 1.640 1.975 2.020 ;
        RECT  1.600 0.550 1.975 0.710 ;
        RECT  2.825 0.550 3.460 0.710 ;
        RECT  2.825 1.640 3.090 2.020 ;
    END
END CKBD6

MACRO CKBD8
    CLASS CORE ;
    FOREIGN CKBD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.265 ;
        END
    END CLK
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.650 2.510 2.030 ;
        RECT  1.660 0.470 2.510 0.630 ;
        RECT  2.510 0.470 2.930 2.030 ;
        RECT  2.930 1.650 3.570 2.030 ;
        RECT  2.930 0.470 3.580 0.630 ;
        RECT  3.570 1.870 4.420 2.030 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.430 0.300 ;
        RECT  0.430 -0.300 0.650 0.340 ;
        RECT  0.650 -0.300 1.270 0.300 ;
        RECT  1.270 -0.300 1.490 0.340 ;
        RECT  1.490 -0.300 2.100 0.300 ;
        RECT  2.100 -0.300 2.320 0.340 ;
        RECT  2.320 -0.300 2.930 0.300 ;
        RECT  2.930 -0.300 3.150 0.340 ;
        RECT  3.150 -0.300 3.750 0.300 ;
        RECT  3.750 -0.300 3.970 0.340 ;
        RECT  3.970 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.290 2.820 ;
        RECT  1.290 2.180 1.510 2.820 ;
        RECT  1.510 2.220 2.110 2.820 ;
        RECT  2.110 2.180 2.330 2.820 ;
        RECT  2.330 2.220 2.930 2.820 ;
        RECT  2.930 2.180 3.150 2.820 ;
        RECT  3.150 2.220 3.760 2.820 ;
        RECT  3.760 2.180 3.980 2.820 ;
        RECT  3.980 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.070 0.885 2.190 1.045 ;
        RECT  1.070 1.960 1.100 2.100 ;
        RECT  1.040 0.885 1.070 2.100 ;
        RECT  0.910 0.440 1.040 2.100 ;
        RECT  0.880 0.440 0.910 1.045 ;
        RECT  0.250 1.390 0.910 1.510 ;
        RECT  0.880 1.960 0.910 2.100 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.090 1.390 0.250 2.100 ;
        RECT  0.060 1.960 0.090 2.100 ;
        LAYER M1 ;
        RECT  3.570 1.870 4.420 2.030 ;
        RECT  1.660 0.470 2.295 0.630 ;
        RECT  1.700 1.650 2.295 2.030 ;
        RECT  3.145 0.470 3.580 0.630 ;
        RECT  3.145 1.650 3.570 2.030 ;
    END
END CKBD8

MACRO CKLNQD1
    CLASS CORE ;
    FOREIGN CKLNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.960 4.550 2.100 ;
        RECT  4.550 0.660 4.710 2.100 ;
        RECT  4.710 1.960 4.740 2.100 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.005 3.440 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.180 0.300 ;
        RECT  4.180 -0.300 4.400 0.340 ;
        RECT  4.400 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  3.940 0.470 4.100 1.570 ;
        RECT  2.420 0.470 3.940 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  4.400 1.030 4.430 1.270 ;
        RECT  4.250 1.030 4.400 1.850 ;
        RECT  4.000 1.690 4.250 1.850 ;
        RECT  3.780 1.690 4.000 2.100 ;
        RECT  3.720 1.690 3.780 1.850 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  3.560 0.710 3.720 1.850 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
    END
END CKLNQD1

MACRO CKLNQD12
    CLASS CORE ;
    FOREIGN CKLNQD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.190 1.640 6.990 2.020 ;
        RECT  5.190 0.740 6.990 0.900 ;
        RECT  6.990 0.740 7.410 2.020 ;
        RECT  7.410 1.640 8.860 2.020 ;
        RECT  7.410 0.740 8.880 0.900 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.480 ;
        RECT  3.750 1.360 4.650 1.480 ;
        RECT  4.650 1.030 4.810 1.480 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 3.530 0.300 ;
        RECT  3.530 -0.300 3.750 0.340 ;
        RECT  3.750 -0.300 4.790 0.300 ;
        RECT  4.790 -0.300 5.010 0.340 ;
        RECT  5.010 -0.300 5.480 0.300 ;
        RECT  5.480 -0.300 5.700 0.340 ;
        RECT  5.700 -0.300 6.170 0.300 ;
        RECT  6.170 -0.300 6.390 0.340 ;
        RECT  6.390 -0.300 6.860 0.300 ;
        RECT  6.860 -0.300 7.080 0.340 ;
        RECT  7.080 -0.300 7.550 0.300 ;
        RECT  7.550 -0.300 7.770 0.340 ;
        RECT  7.770 -0.300 8.240 0.300 ;
        RECT  8.240 -0.300 8.460 0.340 ;
        RECT  8.460 -0.300 8.930 0.300 ;
        RECT  8.930 -0.300 9.150 0.340 ;
        RECT  9.150 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  4.000 1.080 4.230 1.240 ;
        RECT  3.880 0.470 4.000 1.240 ;
        RECT  2.420 0.470 3.880 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  5.060 1.080 6.380 1.240 ;
        RECT  4.940 0.710 5.060 1.780 ;
        RECT  4.120 0.710 4.940 0.870 ;
        RECT  4.720 1.640 4.940 1.780 ;
        RECT  4.500 1.640 4.720 2.060 ;
        RECT  4.030 1.640 4.500 1.780 ;
        RECT  3.810 1.640 4.030 2.060 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        LAYER M1 ;
        RECT  5.190 0.740 6.775 0.900 ;
        RECT  5.190 1.640 6.775 2.020 ;
        RECT  7.625 0.740 8.880 0.900 ;
        RECT  7.625 1.640 8.860 2.020 ;
    END
END CKLNQD12

MACRO CKLNQD16
    CLASS CORE ;
    FOREIGN CKLNQD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.640 8.590 2.020 ;
        RECT  6.050 0.480 8.590 0.640 ;
        RECT  8.590 0.480 9.010 2.020 ;
        RECT  9.010 1.640 11.100 2.020 ;
        RECT  9.010 0.480 11.120 0.640 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.355 3.290 1.515 ;
        RECT  3.290 1.285 3.750 1.515 ;
        RECT  3.750 1.390 4.390 1.510 ;
        RECT  4.390 1.050 4.550 1.510 ;
        RECT  4.550 1.390 5.530 1.510 ;
        RECT  5.530 1.030 5.690 1.510 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.340 ;
        RECT  4.580 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 11.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 3.540 2.820 ;
        RECT  3.540 2.180 3.760 2.820 ;
        RECT  3.760 2.220 11.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 1.840 3.410 2.000 ;
        RECT  2.890 0.710 3.390 0.870 ;
        RECT  5.020 0.810 5.180 1.270 ;
        RECT  4.020 0.810 5.020 0.930 ;
        RECT  3.860 0.810 4.020 1.235 ;
        RECT  3.630 0.810 3.860 0.930 ;
        RECT  3.510 0.470 3.630 0.930 ;
        RECT  2.420 0.470 3.510 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  5.930 1.080 7.595 1.240 ;
        RECT  5.810 0.550 5.930 1.780 ;
        RECT  5.240 0.550 5.810 0.690 ;
        RECT  5.550 1.640 5.810 1.780 ;
        RECT  5.330 1.640 5.550 2.060 ;
        RECT  4.860 1.640 5.330 1.780 ;
        RECT  5.020 0.530 5.240 0.690 ;
        RECT  3.890 0.550 5.020 0.690 ;
        RECT  4.640 1.640 4.860 2.060 ;
        RECT  4.170 1.640 4.640 1.780 ;
        RECT  3.950 1.640 4.170 2.060 ;
        RECT  3.750 0.450 3.890 0.690 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        LAYER M1 ;
        RECT  6.050 0.480 8.375 0.640 ;
        RECT  6.050 1.640 8.375 2.020 ;
        RECT  9.225 0.480 11.120 0.640 ;
        RECT  9.225 1.640 11.100 2.020 ;
    END
END CKLNQD16

MACRO CKLNQD2
    CLASS CORE ;
    FOREIGN CKLNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.470 1.960 4.500 2.100 ;
        RECT  4.500 1.390 4.560 2.100 ;
        RECT  4.450 0.710 4.560 0.870 ;
        RECT  4.560 0.710 4.660 2.100 ;
        RECT  4.660 1.960 4.690 2.100 ;
        RECT  4.660 0.710 4.720 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.005 3.440 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.180 0.300 ;
        RECT  4.180 -0.300 4.400 0.340 ;
        RECT  4.400 -0.300 4.770 0.300 ;
        RECT  4.770 -0.300 4.990 0.340 ;
        RECT  4.990 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  3.940 0.470 4.100 1.570 ;
        RECT  2.420 0.470 3.940 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  4.340 1.050 4.440 1.270 ;
        RECT  4.220 1.050 4.340 1.850 ;
        RECT  4.000 1.690 4.220 1.850 ;
        RECT  3.780 1.690 4.000 2.100 ;
        RECT  3.720 1.690 3.780 1.850 ;
        RECT  3.560 0.710 3.720 1.850 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
    END
END CKLNQD2

MACRO CKLNQD20
    CLASS CORE ;
    FOREIGN CKLNQD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.590 1.640 9.550 2.020 ;
        RECT  6.590 0.470 9.550 0.630 ;
        RECT  9.550 0.470 9.970 2.020 ;
        RECT  9.970 1.640 13.020 2.020 ;
        RECT  9.970 0.470 13.040 0.630 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.510 ;
        RECT  3.750 1.390 4.820 1.510 ;
        RECT  4.820 1.030 4.980 1.510 ;
        RECT  4.980 1.390 6.060 1.510 ;
        RECT  6.060 1.030 6.220 1.510 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.800 0.300 ;
        RECT  4.800 -0.300 5.020 0.340 ;
        RECT  5.020 -0.300 6.190 0.300 ;
        RECT  6.190 -0.300 6.410 0.340 ;
        RECT  6.410 -0.300 13.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 13.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  5.460 0.780 5.620 1.270 ;
        RECT  4.340 0.780 5.460 0.900 ;
        RECT  4.180 0.780 4.340 1.270 ;
        RECT  3.990 0.780 4.180 0.900 ;
        RECT  3.870 0.470 3.990 0.900 ;
        RECT  2.420 0.470 3.870 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  6.460 1.080 8.450 1.240 ;
        RECT  6.340 0.470 6.460 1.780 ;
        RECT  4.110 0.470 6.340 0.630 ;
        RECT  6.120 1.640 6.340 1.780 ;
        RECT  5.900 1.640 6.120 2.060 ;
        RECT  5.410 1.640 5.900 1.780 ;
        RECT  5.190 1.640 5.410 2.060 ;
        RECT  4.720 1.640 5.190 1.780 ;
        RECT  4.500 1.640 4.720 2.060 ;
        RECT  4.030 1.640 4.500 1.780 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        RECT  3.810 1.640 4.030 2.060 ;
        LAYER M1 ;
        RECT  6.590 0.470 9.335 0.630 ;
        RECT  6.590 1.640 9.335 2.020 ;
        RECT  10.185 0.470 13.040 0.630 ;
        RECT  10.185 1.640 13.020 2.020 ;
    END
END CKLNQD20

MACRO CKLNQD24
    CLASS CORE ;
    FOREIGN CKLNQD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.640 10.190 2.020 ;
        RECT  6.490 0.470 10.190 0.630 ;
        RECT  10.190 0.470 10.610 2.020 ;
        RECT  10.610 1.640 14.300 2.020 ;
        RECT  10.610 0.470 14.320 0.630 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.510 ;
        RECT  3.750 1.390 4.880 1.510 ;
        RECT  4.880 1.030 5.040 1.510 ;
        RECT  5.040 1.390 5.990 1.510 ;
        RECT  5.990 1.030 6.130 1.510 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.340 ;
        RECT  5.000 -0.300 14.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 14.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.320 2.000 ;
        RECT  5.520 0.780 5.680 1.270 ;
        RECT  4.400 0.780 5.520 0.900 ;
        RECT  4.240 0.780 4.400 1.270 ;
        RECT  3.990 0.780 4.240 0.900 ;
        RECT  3.870 0.470 3.990 0.900 ;
        RECT  2.420 0.470 3.870 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  6.370 1.080 9.310 1.240 ;
        RECT  6.250 0.470 6.370 1.780 ;
        RECT  4.110 0.470 6.250 0.630 ;
        RECT  6.010 1.640 6.250 1.780 ;
        RECT  5.790 1.640 6.010 2.060 ;
        RECT  5.320 1.640 5.790 1.780 ;
        RECT  5.100 1.640 5.320 2.060 ;
        RECT  4.630 1.640 5.100 1.780 ;
        RECT  4.410 1.640 4.630 2.060 ;
        RECT  3.940 1.640 4.410 1.780 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        RECT  3.720 1.640 3.940 2.060 ;
        LAYER M1 ;
        RECT  6.490 0.470 9.975 0.630 ;
        RECT  6.490 1.640 9.975 2.020 ;
        RECT  10.825 0.470 14.320 0.630 ;
        RECT  10.825 1.640 14.300 2.020 ;
    END
END CKLNQD24

MACRO CKLNQD3
    CLASS CORE ;
    FOREIGN CKLNQD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.460 1.640 4.750 2.020 ;
        RECT  4.440 0.740 4.750 0.900 ;
        RECT  4.750 0.740 5.170 2.020 ;
        RECT  5.170 1.640 5.370 2.020 ;
        RECT  5.170 0.740 5.370 0.900 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.005 3.430 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.170 0.300 ;
        RECT  4.170 -0.300 4.390 0.340 ;
        RECT  4.390 -0.300 4.860 0.300 ;
        RECT  4.860 -0.300 5.080 0.340 ;
        RECT  5.080 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  3.930 0.470 4.090 1.510 ;
        RECT  2.420 0.470 3.930 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  4.330 1.080 4.535 1.240 ;
        RECT  4.210 1.080 4.330 1.790 ;
        RECT  3.990 1.650 4.210 1.790 ;
        RECT  3.770 1.650 3.990 2.080 ;
        RECT  3.710 1.650 3.770 1.790 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        RECT  3.550 0.710 3.710 1.790 ;
        LAYER M1 ;
        RECT  4.440 0.740 4.535 0.900 ;
        RECT  4.460 1.640 4.535 2.020 ;
    END
END CKLNQD3

MACRO CKLNQD4
    CLASS CORE ;
    FOREIGN CKLNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.640 5.070 2.020 ;
        RECT  4.530 0.740 5.070 0.900 ;
        RECT  5.070 0.740 5.490 2.020 ;
        RECT  5.490 1.640 5.560 2.020 ;
        RECT  5.490 0.740 5.580 0.900 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 1.005 3.430 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 4.160 0.300 ;
        RECT  4.160 -0.300 4.380 0.340 ;
        RECT  4.380 -0.300 4.950 0.300 ;
        RECT  4.950 -0.300 5.170 0.340 ;
        RECT  5.170 -0.300 5.730 0.300 ;
        RECT  5.730 -0.300 5.950 0.340 ;
        RECT  5.950 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 4.150 2.820 ;
        RECT  4.150 2.180 4.370 2.820 ;
        RECT  4.370 2.220 4.950 2.820 ;
        RECT  4.950 2.180 5.170 2.820 ;
        RECT  5.170 2.220 5.730 2.820 ;
        RECT  5.730 2.180 5.950 2.820 ;
        RECT  5.950 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.600 0.720 2.630 1.850 ;
        RECT  2.510 0.720 2.600 2.100 ;
        RECT  2.440 1.730 2.510 2.100 ;
        RECT  1.540 1.730 2.440 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.340 2.000 ;
        RECT  3.930 0.470 4.090 1.510 ;
        RECT  2.420 0.470 3.930 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  4.330 1.080 4.660 1.240 ;
        RECT  4.210 1.080 4.330 1.790 ;
        RECT  3.960 1.650 4.210 1.790 ;
        RECT  3.740 1.650 3.960 2.080 ;
        RECT  3.710 1.650 3.740 1.790 ;
        RECT  3.550 0.710 3.710 1.790 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        LAYER M1 ;
        RECT  4.530 0.740 4.855 0.900 ;
        RECT  4.550 1.640 4.855 2.020 ;
    END
END CKLNQD4

MACRO CKLNQD6
    CLASS CORE ;
    FOREIGN CKLNQD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.640 6.030 2.020 ;
        RECT  5.280 0.740 6.030 0.900 ;
        RECT  6.030 0.740 6.450 2.020 ;
        RECT  6.450 1.640 6.920 2.020 ;
        RECT  6.450 0.740 6.940 0.900 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.480 ;
        RECT  3.750 1.360 4.760 1.480 ;
        RECT  4.760 1.030 4.920 1.480 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 3.570 0.300 ;
        RECT  3.570 -0.300 3.790 0.340 ;
        RECT  3.790 -0.300 4.880 0.300 ;
        RECT  4.880 -0.300 5.100 0.340 ;
        RECT  5.100 -0.300 5.590 0.300 ;
        RECT  5.590 -0.300 5.810 0.340 ;
        RECT  5.810 -0.300 6.300 0.300 ;
        RECT  6.300 -0.300 6.520 0.340 ;
        RECT  6.520 -0.300 7.010 0.300 ;
        RECT  7.010 -0.300 7.230 0.340 ;
        RECT  7.230 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 3.470 2.820 ;
        RECT  3.470 2.180 3.690 2.820 ;
        RECT  3.690 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  4.060 1.080 4.340 1.240 ;
        RECT  3.940 0.470 4.060 1.240 ;
        RECT  2.420 0.470 3.940 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  5.160 1.080 5.770 1.240 ;
        RECT  5.040 0.710 5.160 1.780 ;
        RECT  4.210 0.710 5.040 0.870 ;
        RECT  4.780 1.640 5.040 1.780 ;
        RECT  4.560 1.640 4.780 2.060 ;
        RECT  4.090 1.640 4.560 1.780 ;
        RECT  3.870 1.640 4.090 2.060 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        LAYER M1 ;
        RECT  6.665 1.640 6.920 2.020 ;
        RECT  5.280 1.640 5.815 2.020 ;
        RECT  6.665 0.740 6.940 0.900 ;
        RECT  5.280 0.740 5.815 0.900 ;
    END
END CKLNQD6

MACRO CKLNQD8
    CLASS CORE ;
    FOREIGN CKLNQD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.930 0.550 1.515 ;
        RECT  0.550 0.930 0.760 1.090 ;
        END
    END TE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.640 6.350 2.020 ;
        RECT  5.280 0.740 6.350 0.900 ;
        RECT  6.350 0.740 6.770 2.020 ;
        RECT  6.770 1.640 7.580 2.020 ;
        RECT  6.770 0.740 7.600 0.900 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END E
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.480 ;
        RECT  3.750 1.360 4.760 1.480 ;
        RECT  4.760 1.030 4.920 1.480 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.340 ;
        RECT  2.990 -0.300 3.540 0.300 ;
        RECT  3.540 -0.300 3.760 0.340 ;
        RECT  3.760 -0.300 4.880 0.300 ;
        RECT  4.880 -0.300 5.100 0.340 ;
        RECT  5.100 -0.300 5.580 0.300 ;
        RECT  5.580 -0.300 5.800 0.340 ;
        RECT  5.800 -0.300 6.270 0.300 ;
        RECT  6.270 -0.300 6.490 0.340 ;
        RECT  6.490 -0.300 6.960 0.300 ;
        RECT  6.960 -0.300 7.180 0.340 ;
        RECT  7.180 -0.300 7.650 0.300 ;
        RECT  7.650 -0.300 7.870 0.340 ;
        RECT  7.870 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.730 2.820 ;
        RECT  1.730 1.970 1.950 2.820 ;
        RECT  1.950 2.220 3.480 2.820 ;
        RECT  3.480 2.180 3.700 2.820 ;
        RECT  3.700 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.000 ;
        RECT  1.910 0.710 2.010 0.830 ;
        RECT  1.790 0.480 1.910 0.830 ;
        RECT  1.290 0.480 1.790 0.640 ;
        RECT  1.170 0.480 1.290 1.610 ;
        RECT  1.140 0.480 1.170 0.640 ;
        RECT  2.510 0.720 2.630 2.050 ;
        RECT  2.290 1.890 2.510 2.050 ;
        RECT  2.170 1.730 2.290 2.050 ;
        RECT  1.540 1.730 2.170 1.850 ;
        RECT  1.540 0.760 1.660 0.920 ;
        RECT  1.420 0.760 1.540 1.850 ;
        RECT  0.890 1.730 1.420 1.850 ;
        RECT  0.890 1.110 1.050 1.330 ;
        RECT  2.890 0.710 3.410 0.870 ;
        RECT  2.890 1.840 3.350 2.000 ;
        RECT  4.070 1.080 4.300 1.240 ;
        RECT  3.950 0.470 4.070 1.240 ;
        RECT  2.420 0.470 3.950 0.590 ;
        RECT  2.390 0.420 2.420 0.590 ;
        RECT  2.320 0.420 2.390 1.260 ;
        RECT  2.270 0.420 2.320 1.610 ;
        RECT  2.180 0.420 2.270 0.590 ;
        RECT  2.160 1.120 2.270 1.610 ;
        RECT  5.160 1.080 6.085 1.240 ;
        RECT  5.040 0.730 5.160 1.780 ;
        RECT  4.210 0.730 5.040 0.890 ;
        RECT  4.800 1.640 5.040 1.780 ;
        RECT  4.580 1.640 4.800 2.060 ;
        RECT  4.100 1.640 4.580 1.780 ;
        RECT  3.880 1.640 4.100 2.060 ;
        RECT  1.660 1.120 2.160 1.280 ;
        RECT  2.750 0.710 2.890 2.000 ;
        RECT  0.770 1.210 0.890 1.850 ;
        RECT  1.010 1.450 1.170 1.610 ;
        RECT  0.070 0.490 1.000 0.645 ;
        LAYER M1 ;
        RECT  6.985 1.640 7.580 2.020 ;
        RECT  6.985 0.740 7.600 0.900 ;
        RECT  5.280 1.640 6.135 2.020 ;
        RECT  5.280 0.740 6.135 0.900 ;
    END
END CKLNQD8

MACRO CKMUX2D0
    CLASS CORE ;
    FOREIGN CKMUX2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.660 2.790 2.100 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.640 ;
        RECT  0.760 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.940 0.670 2.820 ;
        RECT  0.670 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.890 0.710 2.000 0.870 ;
        RECT  1.890 1.650 2.020 1.810 ;
        RECT  0.060 1.660 0.380 1.820 ;
        RECT  0.350 0.760 0.380 0.880 ;
        RECT  0.380 0.760 0.500 1.820 ;
        RECT  0.500 1.700 0.790 1.820 ;
        RECT  0.790 1.700 0.910 2.050 ;
        RECT  0.910 1.930 1.560 2.050 ;
        RECT  1.560 1.930 1.800 2.100 ;
        RECT  1.030 0.590 1.190 1.760 ;
        RECT  2.460 1.050 2.510 1.290 ;
        RECT  2.340 0.470 2.460 1.290 ;
        RECT  1.570 0.470 2.340 0.590 ;
        RECT  1.410 0.470 1.570 1.760 ;
        RECT  1.760 0.710 1.890 1.810 ;
        RECT  0.190 0.430 0.350 0.880 ;
        RECT  0.920 0.590 1.030 0.750 ;
        RECT  1.320 0.470 1.410 0.630 ;
    END
END CKMUX2D0

MACRO CKMUX2D1
    CLASS CORE ;
    FOREIGN CKMUX2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.610 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.640 ;
        RECT  0.760 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.970 0.670 2.820 ;
        RECT  0.670 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.410 0.470 1.570 1.760 ;
        RECT  1.570 0.470 2.340 0.590 ;
        RECT  2.340 0.470 2.460 1.290 ;
        RECT  2.460 1.050 2.510 1.290 ;
        RECT  1.890 0.710 2.000 0.870 ;
        RECT  1.890 1.640 2.020 1.800 ;
        RECT  0.060 1.690 0.380 1.850 ;
        RECT  0.350 0.760 0.380 0.880 ;
        RECT  0.380 0.760 0.500 1.850 ;
        RECT  0.500 1.730 0.790 1.850 ;
        RECT  0.790 1.730 0.910 2.050 ;
        RECT  0.910 1.930 1.560 2.050 ;
        RECT  1.560 1.930 1.800 2.100 ;
        RECT  1.030 0.590 1.190 1.760 ;
        RECT  1.320 0.470 1.410 0.630 ;
        RECT  1.760 0.710 1.890 1.800 ;
        RECT  0.190 0.430 0.350 0.880 ;
        RECT  0.920 0.590 1.030 0.750 ;
    END
END CKMUX2D1

MACRO CKMUX2D2
    CLASS CORE ;
    FOREIGN CKMUX2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.960 2.550 2.100 ;
        RECT  2.550 1.390 2.650 2.100 ;
        RECT  2.550 0.660 2.650 0.910 ;
        RECT  2.650 0.660 2.710 2.100 ;
        RECT  2.710 1.960 2.740 2.100 ;
        RECT  2.710 0.790 2.790 1.515 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.640 ;
        RECT  0.760 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.940 0.670 2.820 ;
        RECT  0.670 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.910 1.930 1.560 2.050 ;
        RECT  1.560 1.930 1.800 2.100 ;
        RECT  1.030 0.590 1.190 1.760 ;
        RECT  0.790 1.700 0.910 2.050 ;
        RECT  0.500 1.700 0.790 1.820 ;
        RECT  0.380 0.760 0.500 1.820 ;
        RECT  0.350 0.760 0.380 0.880 ;
        RECT  0.060 1.660 0.380 1.820 ;
        RECT  1.890 1.640 2.020 1.800 ;
        RECT  1.890 0.710 2.000 0.870 ;
        RECT  2.430 1.080 2.530 1.240 ;
        RECT  2.310 0.470 2.430 1.240 ;
        RECT  1.570 0.470 2.310 0.590 ;
        RECT  1.410 0.470 1.570 1.760 ;
        RECT  1.320 0.470 1.410 0.630 ;
        RECT  1.760 0.710 1.890 1.800 ;
        RECT  0.190 0.440 0.350 0.880 ;
        RECT  0.920 0.590 1.030 0.750 ;
    END
END CKMUX2D2

MACRO CKMUX2D4
    CLASS CORE ;
    FOREIGN CKMUX2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.650 3.790 2.030 ;
        RECT  3.470 0.690 3.790 0.850 ;
        RECT  3.790 0.690 4.210 2.030 ;
        RECT  4.210 1.650 4.380 2.030 ;
        RECT  4.210 0.690 4.400 0.850 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.005 2.480 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.005 3.110 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.560 0.300 ;
        RECT  0.560 -0.300 0.780 0.340 ;
        RECT  0.780 -0.300 2.490 0.300 ;
        RECT  2.490 -0.300 2.710 0.340 ;
        RECT  2.710 -0.300 3.180 0.300 ;
        RECT  3.180 -0.300 3.400 0.340 ;
        RECT  3.400 -0.300 3.760 0.300 ;
        RECT  3.760 -0.300 3.980 0.340 ;
        RECT  3.980 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.260 0.720 1.190 0.880 ;
        RECT  0.900 1.390 1.060 1.930 ;
        RECT  0.260 1.390 0.900 1.510 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.140 0.720 0.260 2.100 ;
        RECT  0.100 1.390 0.140 2.100 ;
        RECT  2.200 1.650 2.330 1.810 ;
        RECT  2.200 0.710 2.320 0.870 ;
        RECT  2.080 0.710 2.200 1.810 ;
        RECT  2.810 0.710 3.020 0.870 ;
        RECT  2.810 1.890 3.020 2.050 ;
        RECT  2.690 0.710 2.810 2.050 ;
        RECT  1.860 1.930 2.690 2.050 ;
        RECT  1.810 0.720 1.950 0.880 ;
        RECT  1.810 1.430 1.860 2.050 ;
        RECT  1.700 0.720 1.810 2.050 ;
        RECT  3.350 1.080 3.575 1.240 ;
        RECT  3.230 0.470 3.350 1.240 ;
        RECT  1.570 0.470 3.230 0.590 ;
        RECT  1.480 0.470 1.570 0.880 ;
        RECT  1.450 0.470 1.480 1.930 ;
        RECT  1.690 0.720 1.700 1.550 ;
        RECT  1.320 0.720 1.450 1.930 ;
        RECT  1.930 1.100 2.080 1.260 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  3.470 0.690 3.575 0.850 ;
        RECT  3.470 1.650 3.575 2.030 ;
    END
END CKMUX2D4

MACRO CKND0
    CLASS CORE ;
    FOREIGN CKND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.960 0.710 2.100 ;
        RECT  0.710 0.660 0.870 2.100 ;
        RECT  0.870 1.960 0.900 2.100 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.220 0.300 ;
        RECT  0.220 -0.300 0.440 0.340 ;
        RECT  0.440 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.220 2.820 ;
        RECT  0.220 2.180 0.440 2.820 ;
        RECT  0.440 2.220 0.960 2.820 ;
        END
    END VDD
END CKND0

MACRO CKND1
    CLASS CORE ;
    FOREIGN CKND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.960 0.560 2.100 ;
        RECT  0.530 0.435 0.690 0.915 ;
        RECT  0.560 1.390 0.720 2.100 ;
        RECT  0.690 0.795 0.720 0.915 ;
        RECT  0.720 1.960 0.750 2.100 ;
        RECT  0.720 0.795 0.880 1.515 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.290 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.910 0.300 ;
        RECT  0.910 -0.300 1.130 0.340 ;
        RECT  1.130 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.930 2.820 ;
        RECT  0.930 2.180 1.150 2.820 ;
        RECT  1.150 2.220 1.280 2.820 ;
        END
    END VDD
END CKND1

MACRO CKND12
    CLASS CORE ;
    FOREIGN CKND12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.820 0.940 1.980 ;
        RECT  0.940 1.600 3.790 1.980 ;
        RECT  0.720 0.470 3.790 0.690 ;
        RECT  3.790 0.470 4.210 1.980 ;
        RECT  4.210 1.600 6.760 1.980 ;
        RECT  6.760 1.820 7.580 1.980 ;
        RECT  4.210 0.470 7.610 0.690 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.480 0.250 1.235 ;
        RECT  0.250 0.860 2.670 1.020 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 2.180 0.760 2.820 ;
        RECT  0.760 2.220 6.940 2.820 ;
        RECT  6.940 2.180 7.160 2.820 ;
        RECT  7.160 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.760 1.820 7.580 1.980 ;
        RECT  0.940 1.600 3.575 1.980 ;
        RECT  0.720 0.470 3.575 0.690 ;
        RECT  4.425 0.470 7.610 0.690 ;
        RECT  0.120 1.820 0.940 1.980 ;
        RECT  4.425 1.600 6.760 1.980 ;
    END
END CKND12

MACRO CKND16
    CLASS CORE ;
    FOREIGN CKND16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.160 1.600 4.750 1.980 ;
        RECT  0.750 0.470 4.750 0.710 ;
        RECT  4.750 0.470 5.170 1.980 ;
        RECT  5.170 0.470 9.440 0.710 ;
        RECT  5.170 1.600 9.790 1.980 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.480 0.250 1.235 ;
        RECT  0.250 0.880 3.885 1.040 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.560 2.820 ;
        RECT  0.560 2.180 0.780 2.820 ;
        RECT  0.780 2.220 9.170 2.820 ;
        RECT  9.170 2.180 9.390 2.820 ;
        RECT  9.390 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.470 4.535 0.710 ;
        RECT  5.385 0.470 9.440 0.710 ;
        RECT  0.160 1.600 4.535 1.980 ;
        RECT  5.385 1.600 9.790 1.980 ;
    END
END CKND16

MACRO CKND2
    CLASS CORE ;
    FOREIGN CKND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.960 0.510 2.100 ;
        RECT  0.510 1.390 0.670 2.100 ;
        RECT  0.670 1.960 0.700 2.100 ;
        RECT  0.670 1.390 1.040 1.515 ;
        RECT  1.040 0.435 1.200 1.515 ;
        RECT  1.220 1.960 1.250 2.100 ;
        RECT  1.200 1.390 1.250 1.515 ;
        RECT  1.250 1.390 1.410 2.100 ;
        RECT  1.410 1.960 1.440 2.100 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.290 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.600 0.300 ;
        RECT  0.600 -0.300 0.820 0.340 ;
        RECT  0.820 -0.300 1.420 0.300 ;
        RECT  1.420 -0.300 1.640 0.340 ;
        RECT  1.640 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
END CKND2

MACRO CKND20
    CLASS CORE ;
    FOREIGN CKND20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.640 5.710 2.020 ;
        RECT  0.750 0.470 5.710 0.710 ;
        RECT  5.710 0.470 6.130 2.020 ;
        RECT  6.130 1.640 11.620 2.020 ;
        RECT  6.130 0.470 11.680 0.710 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.480 0.230 1.515 ;
        RECT  0.230 0.480 0.250 1.040 ;
        RECT  0.250 0.880 4.885 1.040 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 2.180 0.760 2.820 ;
        RECT  0.760 2.220 11.800 2.820 ;
        RECT  11.800 2.180 12.020 2.820 ;
        RECT  12.020 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 0.470 5.495 0.710 ;
        RECT  6.345 0.470 11.680 0.710 ;
        RECT  0.140 1.640 5.495 2.020 ;
        RECT  6.345 1.640 11.620 2.020 ;
    END
END CKND20

MACRO CKND24
    CLASS CORE ;
    FOREIGN CKND24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.150 1.600 6.670 1.980 ;
        RECT  0.730 0.470 6.670 0.710 ;
        RECT  6.670 0.470 7.090 1.980 ;
        RECT  7.090 1.600 13.860 1.980 ;
        RECT  7.090 0.470 13.920 0.710 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.480 0.230 1.235 ;
        RECT  0.230 0.480 0.250 1.040 ;
        RECT  0.250 0.880 5.885 1.040 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 14.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.550 2.820 ;
        RECT  0.550 2.180 0.770 2.820 ;
        RECT  0.770 2.220 14.040 2.820 ;
        RECT  14.040 2.180 14.260 2.820 ;
        RECT  14.260 2.220 14.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.305 0.470 13.920 0.710 ;
        RECT  0.730 0.470 6.455 0.710 ;
        RECT  0.150 1.600 6.455 1.980 ;
        RECT  7.305 1.600 13.860 1.980 ;
    END
END CKND24

MACRO CKND2D0
    CLASS CORE ;
    FOREIGN CKND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.640 1.050 1.800 ;
        RECT  0.790 0.720 1.050 0.880 ;
        RECT  1.050 0.720 1.190 1.800 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.930 2.820 ;
        RECT  0.930 2.180 1.150 2.820 ;
        RECT  1.150 2.220 1.280 2.820 ;
        END
    END VDD
END CKND2D0

MACRO CKND2D1
    CLASS CORE ;
    FOREIGN CKND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.960 0.560 2.100 ;
        RECT  0.560 1.390 0.720 2.100 ;
        RECT  0.720 1.960 0.750 2.100 ;
        RECT  0.720 1.390 1.050 1.515 ;
        RECT  0.790 0.550 1.050 0.710 ;
        RECT  1.050 0.550 1.190 1.515 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.930 2.820 ;
        RECT  0.930 2.180 1.150 2.820 ;
        RECT  1.150 2.220 1.280 2.820 ;
        END
    END VDD
END CKND2D1

MACRO CKND2D2
    CLASS CORE ;
    FOREIGN CKND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.470 0.550 1.650 ;
        RECT  0.550 0.470 1.190 0.630 ;
        RECT  0.550 1.490 1.450 1.650 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.890 ;
        RECT  0.250 1.770 1.570 1.890 ;
        RECT  1.330 1.060 1.570 1.220 ;
        RECT  1.570 1.060 1.690 1.890 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.190 0.300 ;
        RECT  0.190 -0.300 0.410 0.340 ;
        RECT  0.410 -0.300 1.510 0.300 ;
        RECT  1.510 -0.300 1.730 0.340 ;
        RECT  1.730 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
END CKND2D2

MACRO CKND2D3
    CLASS CORE ;
    FOREIGN CKND2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.600 0.670 2.020 ;
        RECT  0.820 0.450 1.060 0.605 ;
        RECT  0.670 1.600 1.140 1.730 ;
        RECT  1.140 1.600 1.360 2.020 ;
        RECT  1.360 1.600 1.870 1.730 ;
        RECT  1.060 0.470 2.200 0.605 ;
        RECT  1.870 1.425 2.290 1.935 ;
        RECT  2.290 1.425 2.360 1.545 ;
        RECT  2.200 0.450 2.360 0.605 ;
        RECT  2.360 0.450 2.480 1.545 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 0.985 0.520 1.475 ;
        RECT  0.520 1.355 1.050 1.475 ;
        RECT  1.050 1.005 1.170 1.475 ;
        RECT  1.170 1.005 1.510 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.235 ;
        RECT  0.870 0.725 2.080 0.845 ;
        RECT  2.080 0.725 2.240 1.135 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.170 0.300 ;
        RECT  0.170 -0.300 0.390 0.340 ;
        RECT  0.390 -0.300 1.540 0.300 ;
        RECT  1.540 -0.300 1.760 0.340 ;
        RECT  1.760 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.360 0.450 2.480 1.210 ;
        RECT  2.200 0.450 2.360 0.605 ;
        RECT  1.060 0.470 2.200 0.605 ;
        RECT  1.360 1.600 1.655 1.730 ;
        RECT  1.140 1.600 1.360 2.020 ;
        RECT  0.670 1.600 1.140 1.730 ;
        RECT  0.450 1.600 0.670 2.020 ;
        RECT  0.820 0.450 1.060 0.605 ;
    END
END CKND2D3

MACRO CKND2D4
    CLASS CORE ;
    FOREIGN CKND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.960 0.450 2.100 ;
        RECT  0.450 0.710 0.610 2.100 ;
        RECT  0.610 1.880 0.640 2.100 ;
        RECT  0.610 0.710 1.020 0.870 ;
        RECT  0.640 1.880 1.130 2.040 ;
        RECT  1.130 1.630 1.350 2.040 ;
        RECT  1.350 1.880 1.830 2.040 ;
        RECT  1.830 1.630 2.050 2.040 ;
        RECT  2.050 1.880 2.510 2.040 ;
        RECT  2.510 1.425 2.650 2.040 ;
        RECT  2.150 0.730 2.650 0.890 ;
        RECT  2.650 0.730 2.790 2.040 ;
        RECT  2.790 1.425 2.930 2.040 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.470 0.250 1.290 ;
        RECT  0.250 0.470 1.520 0.590 ;
        RECT  1.520 0.470 1.680 1.270 ;
        RECT  1.680 0.470 2.910 0.590 ;
        RECT  2.910 0.470 3.070 1.250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.030 1.235 ;
        RECT  1.030 1.005 1.190 1.510 ;
        RECT  1.190 1.390 2.010 1.510 ;
        RECT  2.010 1.030 2.170 1.510 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.480 0.300 ;
        RECT  1.480 -0.300 1.700 0.340 ;
        RECT  1.700 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 0.730 2.650 0.890 ;
        RECT  0.420 1.960 0.450 2.100 ;
        RECT  0.450 0.710 0.610 2.100 ;
        RECT  0.610 1.880 0.640 2.100 ;
        RECT  0.610 0.710 1.020 0.870 ;
        RECT  0.640 1.880 1.130 2.040 ;
        RECT  1.130 1.630 1.350 2.040 ;
        RECT  1.350 1.880 1.830 2.040 ;
        RECT  1.830 1.630 2.050 2.040 ;
        RECT  2.050 1.880 2.295 2.040 ;
        RECT  2.650 0.730 2.790 1.210 ;
    END
END CKND2D4

MACRO CKND2D8
    CLASS CORE ;
    FOREIGN CKND2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.600 0.730 1.760 ;
        RECT  0.730 0.480 0.870 1.760 ;
        RECT  0.870 1.600 1.360 1.760 ;
        RECT  1.820 1.570 2.190 1.730 ;
        RECT  2.190 1.145 2.470 1.730 ;
        RECT  0.870 0.480 2.470 0.640 ;
        RECT  2.470 0.480 2.610 1.730 ;
        RECT  2.610 1.570 2.800 1.730 ;
        RECT  3.260 1.600 3.620 1.760 ;
        RECT  2.610 0.765 3.620 0.885 ;
        RECT  3.620 0.765 3.635 1.760 ;
        RECT  3.635 0.480 3.760 1.760 ;
        RECT  3.760 1.600 4.240 1.760 ;
        RECT  4.700 1.600 5.530 1.760 ;
        RECT  3.760 0.480 5.530 0.640 ;
        RECT  5.530 0.480 5.670 1.760 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 2.020 ;
        RECT  0.250 1.900 1.520 2.020 ;
        RECT  1.520 1.030 1.680 2.020 ;
        RECT  1.680 1.900 2.960 2.020 ;
        RECT  2.960 1.005 3.120 2.020 ;
        RECT  3.120 1.900 4.400 2.020 ;
        RECT  4.400 1.050 4.560 2.020 ;
        RECT  4.560 1.900 5.830 2.020 ;
        RECT  5.830 1.005 5.990 2.020 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.880 0.810 4.040 1.290 ;
        RECT  4.040 0.810 4.890 0.930 ;
        RECT  4.890 0.810 5.010 1.235 ;
        RECT  5.010 1.005 5.350 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.450 0.300 ;
        RECT  1.450 -0.300 1.670 0.340 ;
        RECT  1.670 -0.300 2.960 0.300 ;
        RECT  2.960 -0.300 3.180 0.645 ;
        RECT  3.180 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.340 ;
        RECT  4.580 -0.300 5.720 0.300 ;
        RECT  5.720 -0.300 5.940 0.340 ;
        RECT  5.940 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 0.780 2.180 0.960 ;
        RECT  1.150 0.780 1.940 0.900 ;
        RECT  0.990 0.780 1.150 1.290 ;
        LAYER M1 ;
        RECT  3.760 0.480 5.530 0.640 ;
        RECT  5.530 0.480 5.670 1.760 ;
        RECT  4.700 1.600 5.530 1.760 ;
        RECT  3.760 1.600 4.240 1.760 ;
        RECT  3.620 0.480 3.760 1.760 ;
        RECT  2.610 0.765 3.620 0.885 ;
        RECT  3.260 1.600 3.620 1.760 ;
        RECT  2.470 0.480 2.610 0.930 ;
        RECT  0.870 0.480 2.470 0.640 ;
        RECT  0.870 1.600 1.360 1.760 ;
        RECT  0.730 0.480 0.870 1.760 ;
        RECT  1.820 1.570 1.975 1.730 ;
        RECT  0.400 1.600 0.730 1.760 ;
    END
END CKND2D8

MACRO CKND3
    CLASS CORE ;
    FOREIGN CKND3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.640 1.230 2.020 ;
        RECT  0.840 0.500 1.230 0.880 ;
        RECT  1.230 0.500 1.650 2.020 ;
        RECT  1.650 0.500 1.890 0.880 ;
        RECT  1.650 1.640 2.110 2.020 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.290 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.430 0.300 ;
        RECT  0.430 -0.300 0.650 0.340 ;
        RECT  0.650 -0.300 1.260 0.300 ;
        RECT  1.260 -0.300 1.480 0.340 ;
        RECT  1.480 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.865 1.640 2.110 2.020 ;
        RECT  0.450 1.640 1.015 2.020 ;
        RECT  1.865 0.500 1.890 0.880 ;
        RECT  0.840 0.500 1.015 0.880 ;
    END
END CKND3

MACRO CKND4
    CLASS CORE ;
    FOREIGN CKND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 1.230 2.020 ;
        RECT  0.840 0.500 1.230 0.880 ;
        RECT  1.230 0.500 1.650 2.020 ;
        RECT  1.650 0.500 1.890 0.880 ;
        RECT  1.650 1.640 2.760 2.020 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.250 1.290 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.430 0.300 ;
        RECT  0.430 -0.300 0.650 0.340 ;
        RECT  0.650 -0.300 1.260 0.300 ;
        RECT  1.260 -0.300 1.480 0.340 ;
        RECT  1.480 -0.300 2.080 0.300 ;
        RECT  2.080 -0.300 2.300 0.340 ;
        RECT  2.300 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.865 0.500 1.890 0.880 ;
        RECT  0.440 1.640 1.015 2.020 ;
        RECT  1.865 1.640 2.760 2.020 ;
        RECT  0.840 0.500 1.015 0.880 ;
    END
END CKND4

MACRO CKND6
    CLASS CORE ;
    FOREIGN CKND6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.600 1.870 1.980 ;
        RECT  0.860 0.480 1.870 0.860 ;
        RECT  1.870 0.480 2.290 1.980 ;
        RECT  2.290 0.480 2.740 0.860 ;
        RECT  2.290 1.600 4.330 1.980 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.670 0.230 1.515 ;
        RECT  0.230 0.670 0.250 1.240 ;
        RECT  0.250 1.080 1.580 1.240 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 1.280 0.300 ;
        RECT  1.280 -0.300 1.500 0.340 ;
        RECT  1.500 -0.300 2.100 0.300 ;
        RECT  2.100 -0.300 2.320 0.340 ;
        RECT  2.320 -0.300 2.930 0.300 ;
        RECT  2.930 -0.300 3.150 0.340 ;
        RECT  3.150 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.505 1.600 4.330 1.980 ;
        RECT  2.505 0.480 2.740 0.860 ;
        RECT  0.460 1.600 1.655 1.980 ;
        RECT  0.860 0.480 1.655 0.860 ;
    END
END CKND6

MACRO CKND8
    CLASS CORE ;
    FOREIGN CKND8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.960 1.600 2.510 1.980 ;
        RECT  0.810 0.480 2.510 0.640 ;
        RECT  2.510 0.480 2.930 1.980 ;
        RECT  2.930 1.600 5.080 1.980 ;
        RECT  5.080 1.820 5.880 1.980 ;
        RECT  2.930 0.480 5.980 0.640 ;
        END
    END CN
    PIN CLK
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.480 0.230 1.235 ;
        RECT  0.230 0.480 0.250 1.010 ;
        RECT  0.250 0.850 2.225 1.010 ;
        END
    END CLK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.420 0.300 ;
        RECT  0.420 -0.300 0.640 0.340 ;
        RECT  0.640 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 2.080 0.300 ;
        RECT  2.080 -0.300 2.300 0.340 ;
        RECT  2.300 -0.300 2.900 0.300 ;
        RECT  2.900 -0.300 3.120 0.340 ;
        RECT  3.120 -0.300 3.730 0.300 ;
        RECT  3.730 -0.300 3.950 0.340 ;
        RECT  3.950 -0.300 4.540 0.300 ;
        RECT  4.540 -0.300 4.760 0.340 ;
        RECT  4.760 -0.300 5.340 0.300 ;
        RECT  5.340 -0.300 5.560 0.340 ;
        RECT  5.560 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.560 2.820 ;
        RECT  0.560 2.180 0.780 2.820 ;
        RECT  0.780 2.220 1.350 2.820 ;
        RECT  1.350 2.180 1.570 2.820 ;
        RECT  1.570 2.220 2.130 2.820 ;
        RECT  2.130 2.180 2.350 2.820 ;
        RECT  2.350 2.220 2.910 2.820 ;
        RECT  2.910 2.180 3.130 2.820 ;
        RECT  3.130 2.220 3.690 2.820 ;
        RECT  3.690 2.180 3.910 2.820 ;
        RECT  3.910 2.220 4.470 2.820 ;
        RECT  4.470 2.180 4.690 2.820 ;
        RECT  4.690 2.220 5.250 2.820 ;
        RECT  5.250 2.180 5.470 2.820 ;
        RECT  5.470 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.080 1.820 5.880 1.980 ;
        RECT  3.145 0.480 5.980 0.640 ;
        RECT  0.960 1.600 2.295 1.980 ;
        RECT  3.145 1.600 5.080 1.980 ;
        RECT  0.810 0.480 2.295 0.640 ;
    END
END CKND8

MACRO CKXOR2D0
    CLASS CORE ;
    FOREIGN CKXOR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.660 2.790 2.090 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 1.875 0.630 2.820 ;
        RECT  0.630 2.220 2.150 2.820 ;
        RECT  2.150 2.180 2.370 2.820 ;
        RECT  2.370 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.630 0.645 ;
        RECT  0.630 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.750 1.030 0.870 2.050 ;
        RECT  0.870 1.930 1.730 2.050 ;
        RECT  1.730 0.710 1.890 2.050 ;
        RECT  1.890 0.710 2.050 0.870 ;
        RECT  0.100 0.635 0.260 0.885 ;
        RECT  0.260 1.635 0.445 1.755 ;
        RECT  0.260 0.765 0.445 0.885 ;
        RECT  0.445 0.765 0.565 1.755 ;
        RECT  0.565 0.765 0.750 0.885 ;
        RECT  0.750 0.470 0.870 0.885 ;
        RECT  0.870 0.470 1.230 0.590 ;
        RECT  1.230 0.470 1.350 1.385 ;
        RECT  1.110 1.590 1.130 1.810 ;
        RECT  2.350 0.470 2.510 1.345 ;
        RECT  1.610 0.470 2.350 0.590 ;
        RECT  1.300 1.650 1.470 1.810 ;
        RECT  1.470 0.470 1.610 1.810 ;
        RECT  0.710 1.030 0.750 1.270 ;
        RECT  0.100 1.635 0.260 1.875 ;
        RECT  0.990 0.710 1.110 1.810 ;
    END
END CKXOR2D0

MACRO CKXOR2D1
    CLASS CORE ;
    FOREIGN CKXOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.660 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 1.905 0.620 2.820 ;
        RECT  0.620 2.220 2.140 2.820 ;
        RECT  2.140 2.180 2.360 2.820 ;
        RECT  2.360 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.620 0.645 ;
        RECT  0.620 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.350 0.470 2.510 1.290 ;
        RECT  0.740 1.030 0.860 2.050 ;
        RECT  0.860 1.930 1.700 2.050 ;
        RECT  1.700 1.930 1.730 2.100 ;
        RECT  1.730 0.710 1.890 2.100 ;
        RECT  1.890 1.960 1.920 2.100 ;
        RECT  1.890 0.710 2.040 0.870 ;
        RECT  0.090 0.645 0.250 0.885 ;
        RECT  0.250 1.635 0.450 1.755 ;
        RECT  0.250 0.765 0.450 0.885 ;
        RECT  0.450 0.765 0.570 1.755 ;
        RECT  0.570 0.765 0.740 0.885 ;
        RECT  0.740 0.470 0.860 0.885 ;
        RECT  0.860 0.470 1.220 0.590 ;
        RECT  1.220 0.470 1.340 1.290 ;
        RECT  1.100 1.590 1.120 1.810 ;
        RECT  1.600 0.470 2.350 0.590 ;
        RECT  1.460 0.470 1.600 1.810 ;
        RECT  1.290 1.650 1.460 1.810 ;
        RECT  0.720 1.030 0.740 1.270 ;
        RECT  0.090 1.635 0.250 1.880 ;
        RECT  0.980 0.710 1.100 1.810 ;
    END
END CKXOR2D1

MACRO CKXOR2D2
    CLASS CORE ;
    FOREIGN CKXOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.960 2.550 2.100 ;
        RECT  2.550 1.390 2.650 2.100 ;
        RECT  2.550 0.660 2.650 0.900 ;
        RECT  2.650 0.660 2.710 2.100 ;
        RECT  2.710 1.960 2.740 2.100 ;
        RECT  2.710 0.780 2.790 1.515 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 1.905 0.620 2.820 ;
        RECT  0.620 2.220 2.110 2.820 ;
        RECT  2.110 2.180 2.330 2.820 ;
        RECT  2.330 2.220 3.200 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.620 0.645 ;
        RECT  0.620 -0.300 2.120 0.300 ;
        RECT  2.120 -0.300 2.340 0.340 ;
        RECT  2.340 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.200 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.250 0.765 0.450 0.885 ;
        RECT  0.450 0.765 0.570 1.755 ;
        RECT  0.570 0.765 0.740 0.885 ;
        RECT  0.740 0.470 0.860 0.885 ;
        RECT  0.860 0.470 1.220 0.590 ;
        RECT  1.220 0.470 1.340 1.290 ;
        RECT  1.100 1.590 1.120 1.810 ;
        RECT  0.250 1.635 0.450 1.755 ;
        RECT  0.090 0.645 0.250 0.885 ;
        RECT  1.890 0.710 2.040 0.870 ;
        RECT  1.890 1.960 1.920 2.100 ;
        RECT  1.730 0.710 1.890 2.100 ;
        RECT  1.700 1.930 1.730 2.100 ;
        RECT  0.860 1.930 1.700 2.050 ;
        RECT  0.740 1.030 0.860 2.050 ;
        RECT  2.430 1.050 2.490 1.270 ;
        RECT  2.290 0.470 2.430 1.270 ;
        RECT  1.600 0.470 2.290 0.590 ;
        RECT  1.460 0.470 1.600 1.810 ;
        RECT  1.290 1.650 1.460 1.810 ;
        RECT  0.720 1.030 0.740 1.270 ;
        RECT  0.090 1.635 0.250 1.880 ;
        RECT  0.980 0.710 1.100 1.810 ;
    END
END CKXOR2D2

MACRO CKXOR2D4
    CLASS CORE ;
    FOREIGN CKXOR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.650 4.750 2.030 ;
        RECT  4.430 0.710 4.750 0.870 ;
        RECT  4.750 0.710 5.170 2.030 ;
        RECT  5.170 1.650 5.340 2.030 ;
        RECT  5.170 0.710 5.360 0.870 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 4.070 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.485 2.820 ;
        RECT  0.485 2.180 0.705 2.820 ;
        RECT  0.705 2.220 5.760 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 3.230 0.300 ;
        RECT  3.230 -0.300 3.450 0.340 ;
        RECT  3.450 -0.300 4.030 0.300 ;
        RECT  4.030 -0.300 4.250 0.340 ;
        RECT  4.250 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.940 0.340 ;
        RECT  4.940 -0.300 5.410 0.300 ;
        RECT  5.410 -0.300 5.630 0.340 ;
        RECT  5.630 -0.300 5.760 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.110 1.060 1.260 1.280 ;
        RECT  0.990 0.710 1.110 1.800 ;
        RECT  0.840 0.710 0.990 0.870 ;
        RECT  1.760 0.470 1.880 1.560 ;
        RECT  1.660 0.470 1.760 0.635 ;
        RECT  1.620 1.400 1.760 1.560 ;
        RECT  0.260 0.470 1.660 0.590 ;
        RECT  3.770 1.550 3.930 2.050 ;
        RECT  3.420 0.710 3.870 0.870 ;
        RECT  3.420 1.910 3.770 2.050 ;
        RECT  3.300 0.710 3.420 2.050 ;
        RECT  2.570 1.910 3.300 2.050 ;
        RECT  2.570 0.710 2.710 0.870 ;
        RECT  2.410 0.710 2.570 2.050 ;
        RECT  0.520 1.930 2.410 2.050 ;
        RECT  4.310 1.050 4.470 1.270 ;
        RECT  4.190 0.470 4.310 1.270 ;
        RECT  3.040 0.470 4.190 0.590 ;
        RECT  2.880 0.470 3.040 1.710 ;
        RECT  2.290 0.470 2.880 0.590 ;
        RECT  2.740 1.550 2.880 1.710 ;
        RECT  2.170 0.470 2.290 1.810 ;
        RECT  2.050 0.470 2.170 0.630 ;
        RECT  2.000 1.650 2.170 1.810 ;
        RECT  1.500 1.690 2.000 1.810 ;
        RECT  1.380 0.720 1.500 1.810 ;
        RECT  1.240 0.720 1.380 0.940 ;
        RECT  1.240 1.670 1.380 1.810 ;
        RECT  0.380 1.030 0.520 2.050 ;
        RECT  0.100 0.470 0.260 1.960 ;
        RECT  0.860 1.640 0.990 1.800 ;
        LAYER M1 ;
        RECT  4.430 0.710 4.535 0.870 ;
        RECT  4.430 1.650 4.535 2.030 ;
    END
END CKXOR2D4

MACRO CMPE22D1
    CLASS CORE ;
    FOREIGN CMPE22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.180 1.940 4.210 2.100 ;
        RECT  4.210 1.390 4.250 2.100 ;
        RECT  4.210 0.420 4.250 0.920 ;
        RECT  4.250 0.420 4.370 2.100 ;
        RECT  4.370 0.800 4.390 1.515 ;
        RECT  4.370 1.940 4.400 2.100 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 0.440 0.200 2.070 ;
        RECT  0.200 1.565 0.250 2.070 ;
        RECT  0.200 0.440 0.250 0.955 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.080 0.730 1.300 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.360 1.160 1.515 ;
        RECT  1.160 1.360 1.280 2.050 ;
        RECT  1.280 1.930 3.340 2.050 ;
        RECT  3.340 1.930 3.580 2.070 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.080 1.690 1.240 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.220 2.820 ;
        RECT  1.220 2.180 1.440 2.820 ;
        RECT  1.440 2.220 3.780 2.820 ;
        RECT  3.780 2.180 4.000 2.820 ;
        RECT  4.000 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 1.640 2.980 1.810 ;
        RECT  2.850 0.710 2.990 0.850 ;
        RECT  2.980 1.690 3.970 1.810 ;
        RECT  3.970 1.010 4.090 1.810 ;
        RECT  4.090 1.010 4.130 1.230 ;
        RECT  3.490 0.630 3.610 1.560 ;
        RECT  3.610 1.420 3.730 1.560 ;
        RECT  3.610 0.630 3.730 0.790 ;
        RECT  1.670 1.670 2.090 1.810 ;
        RECT  1.920 0.470 2.090 0.590 ;
        RECT  2.090 0.470 2.230 1.810 ;
        RECT  2.230 1.060 2.370 1.280 ;
        RECT  2.230 0.470 3.110 0.590 ;
        RECT  3.110 0.470 3.230 1.540 ;
        RECT  3.230 1.380 3.370 1.540 ;
        RECT  3.230 0.630 3.370 0.790 ;
        RECT  2.370 0.710 2.490 0.850 ;
        RECT  2.490 0.710 2.610 1.810 ;
        RECT  0.370 0.470 0.490 1.785 ;
        RECT  0.490 1.665 0.820 1.785 ;
        RECT  0.820 1.665 1.040 1.825 ;
        RECT  0.490 0.470 1.060 0.590 ;
        RECT  1.060 0.450 1.280 0.870 ;
        RECT  3.350 1.040 3.490 1.200 ;
        RECT  1.700 0.450 1.920 0.870 ;
        RECT  2.730 0.710 2.850 1.810 ;
        RECT  2.360 1.650 2.490 1.810 ;
        RECT  0.320 1.080 0.370 1.300 ;
    END
END CMPE22D1

MACRO CMPE22D2
    CLASS CORE ;
    FOREIGN CMPE22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.760 1.940 4.790 2.100 ;
        RECT  4.790 1.390 4.890 2.100 ;
        RECT  4.790 0.420 4.890 0.900 ;
        RECT  4.890 0.420 4.950 2.100 ;
        RECT  4.950 1.940 4.980 2.100 ;
        RECT  4.950 0.780 5.030 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.805 0.550 1.515 ;
        RECT  0.530 1.940 0.560 2.100 ;
        RECT  0.550 1.390 0.560 1.515 ;
        RECT  0.550 0.805 0.560 0.940 ;
        RECT  0.560 1.390 0.720 2.100 ;
        RECT  0.560 0.440 0.720 0.940 ;
        RECT  0.720 1.940 0.750 2.100 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.080 1.370 1.300 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.360 1.690 1.515 ;
        RECT  1.690 1.360 1.830 2.050 ;
        RECT  1.830 1.930 3.810 2.050 ;
        RECT  3.810 1.930 4.050 2.070 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.080 2.010 1.240 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.080 2.290 1.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.340 ;
        RECT  4.580 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.760 2.820 ;
        RECT  1.760 2.180 1.980 2.820 ;
        RECT  1.980 2.220 4.360 2.820 ;
        RECT  4.360 2.180 4.580 2.820 ;
        RECT  4.580 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.450 1.750 0.870 ;
        RECT  0.960 0.750 1.530 0.870 ;
        RECT  1.290 1.640 1.530 1.800 ;
        RECT  0.960 1.640 1.290 1.760 ;
        RECT  0.840 0.750 0.960 1.760 ;
        RECT  2.960 0.710 3.080 1.810 ;
        RECT  2.840 0.710 2.960 0.850 ;
        RECT  3.700 0.630 3.840 0.790 ;
        RECT  3.700 1.380 3.840 1.540 ;
        RECT  3.580 0.470 3.700 1.540 ;
        RECT  2.700 0.470 3.580 0.590 ;
        RECT  2.700 1.060 2.840 1.280 ;
        RECT  2.560 0.470 2.700 1.810 ;
        RECT  2.390 0.470 2.560 0.590 ;
        RECT  2.140 1.650 2.560 1.810 ;
        RECT  4.080 0.630 4.200 0.790 ;
        RECT  4.080 1.420 4.200 1.560 ;
        RECT  3.960 0.630 4.080 1.560 ;
        RECT  4.670 0.990 4.710 1.230 ;
        RECT  4.550 0.990 4.670 1.810 ;
        RECT  3.450 1.690 4.550 1.810 ;
        RECT  3.320 0.710 3.460 0.850 ;
        RECT  3.320 1.640 3.450 1.810 ;
        RECT  3.200 0.710 3.320 1.810 ;
        RECT  3.820 1.040 3.960 1.200 ;
        RECT  2.170 0.450 2.390 0.870 ;
        RECT  2.830 1.650 2.960 1.810 ;
        RECT  0.720 1.110 0.840 1.270 ;
    END
END CMPE22D2

MACRO CMPE32D1
    CLASS CORE ;
    FOREIGN CMPE32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.680 1.940 7.710 2.100 ;
        RECT  7.710 1.390 7.770 2.100 ;
        RECT  7.710 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.870 2.100 ;
        RECT  7.870 1.940 7.900 2.100 ;
        RECT  7.870 0.780 7.910 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 1.410 7.130 1.550 ;
        RECT  7.010 0.420 7.130 0.900 ;
        RECT  7.130 0.420 7.170 1.550 ;
        RECT  7.170 0.780 7.270 1.550 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 0.725 6.330 1.245 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.040 3.290 1.405 ;
        RECT  3.290 1.285 3.430 1.795 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.940 1.830 4.030 2.050 ;
        RECT  4.000 0.620 4.030 0.860 ;
        RECT  4.030 0.620 4.150 2.050 ;
        RECT  3.650 0.470 3.760 0.690 ;
        RECT  3.760 0.470 3.880 1.630 ;
        RECT  3.880 1.040 3.910 1.260 ;
        RECT  2.260 0.470 2.360 0.630 ;
        RECT  2.260 1.490 2.380 1.650 ;
        RECT  2.360 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.530 1.160 ;
        RECT  3.530 1.020 3.640 1.160 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.830 0.800 1.950 ;
        RECT  0.640 0.760 0.800 0.880 ;
        RECT  0.800 0.760 0.920 1.950 ;
        RECT  0.920 1.090 1.460 1.250 ;
        RECT  0.920 1.830 2.550 1.950 ;
        RECT  2.540 0.710 2.550 0.850 ;
        RECT  2.550 0.710 2.690 1.950 ;
        RECT  2.690 1.470 2.710 1.950 ;
        RECT  2.690 0.710 2.780 0.850 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.090 1.470 1.860 1.630 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.630 ;
        RECT  3.030 1.930 3.940 2.050 ;
        RECT  3.030 0.760 3.150 0.920 ;
        RECT  2.910 0.760 3.030 2.050 ;
        RECT  2.890 1.050 2.910 2.050 ;
        RECT  5.670 0.710 5.800 0.850 ;
        RECT  5.550 0.710 5.670 1.540 ;
        RECT  6.570 0.470 6.690 1.550 ;
        RECT  6.470 0.470 6.570 0.590 ;
        RECT  5.940 1.410 6.570 1.550 ;
        RECT  6.250 0.450 6.470 0.590 ;
        RECT  4.950 0.470 6.250 0.590 ;
        RECT  5.800 1.040 5.940 1.550 ;
        RECT  4.790 0.470 4.950 1.570 ;
        RECT  6.790 1.910 7.030 2.070 ;
        RECT  4.480 1.910 6.790 2.050 ;
        RECT  4.480 0.670 4.590 0.830 ;
        RECT  7.590 1.040 7.650 1.280 ;
        RECT  7.470 1.040 7.590 1.790 ;
        RECT  5.260 1.670 7.470 1.790 ;
        RECT  5.260 0.710 5.400 0.850 ;
        RECT  5.100 0.710 5.260 1.790 ;
        RECT  4.320 0.670 4.480 2.050 ;
        RECT  4.660 1.410 4.790 1.570 ;
        RECT  5.430 1.400 5.550 1.540 ;
        RECT  2.810 1.050 2.890 1.270 ;
        RECT  3.620 1.410 3.760 1.630 ;
        RECT  2.140 0.470 2.260 1.650 ;
        RECT  0.420 1.530 0.640 1.950 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END CMPE32D1

MACRO CMPE32D2
    CLASS CORE ;
    FOREIGN CMPE32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.620 1.940 7.650 2.100 ;
        RECT  7.650 1.390 7.810 2.100 ;
        RECT  7.670 0.420 7.830 0.900 ;
        RECT  7.810 1.940 7.840 2.100 ;
        RECT  7.810 1.390 8.090 1.515 ;
        RECT  7.830 0.780 8.090 0.900 ;
        RECT  8.090 0.780 8.230 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.920 1.940 6.950 2.100 ;
        RECT  6.950 1.390 7.110 2.100 ;
        RECT  7.110 1.390 7.130 1.515 ;
        RECT  6.930 0.745 7.130 0.905 ;
        RECT  7.110 1.940 7.140 2.100 ;
        RECT  7.130 0.745 7.270 1.515 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.330 1.515 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.040 3.290 1.405 ;
        RECT  3.290 1.285 3.430 1.795 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.460 0.710 5.600 1.540 ;
        RECT  5.600 1.400 5.670 1.540 ;
        RECT  5.600 0.710 5.790 0.850 ;
        RECT  2.890 1.050 2.910 2.050 ;
        RECT  2.910 0.760 3.030 2.050 ;
        RECT  3.030 1.480 3.050 2.050 ;
        RECT  3.030 0.760 3.150 0.920 ;
        RECT  3.050 1.930 3.940 2.050 ;
        RECT  3.940 1.830 4.030 2.050 ;
        RECT  4.000 0.620 4.030 0.860 ;
        RECT  4.030 0.620 4.150 2.050 ;
        RECT  3.650 0.640 3.760 0.860 ;
        RECT  3.760 0.640 3.880 1.630 ;
        RECT  3.880 1.040 3.910 1.260 ;
        RECT  2.260 0.470 2.360 0.630 ;
        RECT  2.260 1.490 2.380 1.650 ;
        RECT  2.360 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.530 1.160 ;
        RECT  3.530 1.020 3.640 1.160 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.840 0.800 1.960 ;
        RECT  0.640 0.760 0.800 0.880 ;
        RECT  0.800 0.760 0.920 1.960 ;
        RECT  0.920 1.090 1.460 1.250 ;
        RECT  0.920 1.840 2.540 1.960 ;
        RECT  2.540 0.710 2.680 1.960 ;
        RECT  2.680 1.480 2.710 1.960 ;
        RECT  2.680 0.710 2.780 0.850 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.090 1.470 1.860 1.630 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.630 ;
        RECT  6.030 0.710 6.500 0.870 ;
        RECT  5.940 1.650 6.470 1.810 ;
        RECT  5.940 0.710 6.030 1.170 ;
        RECT  5.910 0.710 5.940 1.810 ;
        RECT  5.800 1.050 5.910 1.810 ;
        RECT  4.900 1.690 5.800 1.810 ;
        RECT  4.900 0.530 4.950 0.770 ;
        RECT  4.780 0.530 4.900 1.810 ;
        RECT  6.800 1.080 6.970 1.240 ;
        RECT  6.680 1.080 6.800 2.050 ;
        RECT  4.480 1.930 6.680 2.050 ;
        RECT  4.480 0.650 4.590 0.810 ;
        RECT  7.550 1.080 7.730 1.240 ;
        RECT  7.430 0.470 7.550 1.240 ;
        RECT  5.330 0.470 7.430 0.590 ;
        RECT  5.310 0.470 5.330 0.820 ;
        RECT  5.190 0.470 5.310 1.570 ;
        RECT  5.050 1.410 5.190 1.570 ;
        RECT  4.320 0.650 4.480 2.050 ;
        RECT  4.660 1.410 4.780 1.570 ;
        RECT  5.450 1.400 5.460 1.540 ;
        RECT  2.810 1.050 2.890 1.270 ;
        RECT  3.620 1.410 3.760 1.630 ;
        RECT  2.140 0.470 2.260 1.650 ;
        RECT  0.420 1.540 0.640 1.960 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END CMPE32D2

MACRO CMPE42D1
    CLASS CORE ;
    FOREIGN CMPE42D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.150 1.940 13.180 2.100 ;
        RECT  13.180 1.390 13.210 2.100 ;
        RECT  13.180 0.420 13.210 0.900 ;
        RECT  13.210 0.420 13.340 2.100 ;
        RECT  13.340 0.780 13.350 1.515 ;
        RECT  13.340 1.940 13.370 2.100 ;
        END
    END S
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.060 9.050 1.405 ;
        RECT  9.050 1.060 9.100 1.795 ;
        RECT  9.100 1.285 9.190 1.795 ;
        END
    END D
    PIN COX
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.870 0.450 7.090 0.870 ;
        RECT  6.870 1.410 7.130 1.550 ;
        RECT  7.090 0.750 7.130 0.870 ;
        RECT  7.130 0.750 7.270 1.550 ;
        END
    END COX
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.420 1.410 12.570 1.550 ;
        RECT  12.420 0.450 12.570 0.870 ;
        RECT  12.570 0.450 12.650 1.550 ;
        RECT  12.650 0.750 12.710 1.550 ;
        END
    END CO
    PIN CIX
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.930 1.005 12.390 1.235 ;
        END
    END CIX
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.005 6.950 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 0.990 2.010 1.210 ;
        RECT  2.010 0.990 2.150 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 0.960 0.300 ;
        RECT  0.960 -0.300 1.180 0.340 ;
        RECT  1.180 -0.300 13.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 0.960 2.820 ;
        RECT  0.960 2.180 1.180 2.820 ;
        RECT  1.180 2.220 13.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.810 1.410 12.280 1.550 ;
        RECT  12.070 0.450 12.290 0.870 ;
        RECT  11.310 0.730 11.430 1.540 ;
        RECT  11.430 1.420 11.520 1.540 ;
        RECT  11.430 0.730 11.550 0.950 ;
        RECT  8.700 1.050 8.720 2.050 ;
        RECT  8.720 0.760 8.840 2.050 ;
        RECT  8.840 0.760 8.960 0.920 ;
        RECT  8.840 1.930 9.770 2.050 ;
        RECT  9.770 1.660 9.890 2.050 ;
        RECT  9.820 0.640 9.890 0.860 ;
        RECT  9.890 0.640 10.010 1.880 ;
        RECT  9.440 0.470 9.570 0.690 ;
        RECT  9.570 0.470 9.600 1.810 ;
        RECT  9.600 0.470 9.690 1.550 ;
        RECT  9.690 1.040 9.770 1.260 ;
        RECT  8.140 0.470 9.100 0.590 ;
        RECT  9.100 0.470 9.220 0.940 ;
        RECT  9.220 0.820 9.320 0.940 ;
        RECT  9.320 0.820 9.440 1.275 ;
        RECT  5.420 0.710 5.430 1.560 ;
        RECT  5.430 0.710 5.550 1.790 ;
        RECT  5.550 0.710 5.660 0.850 ;
        RECT  5.550 1.670 7.300 1.790 ;
        RECT  7.300 1.670 7.420 2.050 ;
        RECT  7.420 1.930 7.440 2.050 ;
        RECT  7.440 1.930 7.660 2.100 ;
        RECT  7.660 1.930 8.350 2.050 ;
        RECT  8.350 0.710 8.490 2.050 ;
        RECT  8.490 1.400 8.520 2.050 ;
        RECT  8.490 0.710 8.590 0.850 ;
        RECT  7.550 0.470 7.710 0.610 ;
        RECT  7.710 0.470 7.830 1.690 ;
        RECT  4.640 0.620 4.660 1.710 ;
        RECT  4.660 0.620 4.800 2.050 ;
        RECT  4.800 1.910 6.680 2.050 ;
        RECT  6.680 1.910 6.920 2.070 ;
        RECT  5.050 0.470 5.210 1.570 ;
        RECT  6.070 1.060 6.170 1.280 ;
        RECT  5.210 0.470 6.170 0.590 ;
        RECT  6.170 0.470 6.310 1.550 ;
        RECT  6.310 0.470 6.520 0.590 ;
        RECT  6.310 1.410 6.730 1.550 ;
        RECT  6.520 0.450 6.740 0.870 ;
        RECT  5.830 0.780 5.950 1.540 ;
        RECT  5.950 0.780 6.050 0.900 ;
        RECT  3.150 1.050 3.170 2.050 ;
        RECT  3.170 0.760 3.310 2.050 ;
        RECT  3.310 0.760 3.410 0.920 ;
        RECT  3.310 1.930 4.220 2.050 ;
        RECT  4.220 1.530 4.290 2.050 ;
        RECT  4.250 0.620 4.290 0.860 ;
        RECT  4.290 0.620 4.340 2.050 ;
        RECT  4.340 0.620 4.410 1.750 ;
        RECT  3.910 0.450 3.970 0.950 ;
        RECT  3.970 0.450 4.050 1.810 ;
        RECT  4.050 0.450 4.090 1.550 ;
        RECT  4.090 1.040 4.170 1.260 ;
        RECT  2.520 0.470 2.620 0.630 ;
        RECT  2.520 1.490 2.640 1.650 ;
        RECT  2.620 0.470 3.670 0.590 ;
        RECT  3.670 0.470 3.790 1.275 ;
        RECT  3.790 1.055 3.850 1.275 ;
        RECT  0.550 0.460 0.770 0.880 ;
        RECT  0.770 1.895 1.070 2.015 ;
        RECT  0.770 0.760 1.070 0.880 ;
        RECT  1.070 0.760 1.190 2.015 ;
        RECT  1.190 1.060 1.320 1.280 ;
        RECT  1.190 1.895 2.800 2.015 ;
        RECT  2.800 0.710 2.940 2.015 ;
        RECT  2.940 1.470 2.970 2.015 ;
        RECT  2.940 0.710 3.040 0.850 ;
        RECT  1.370 0.460 1.490 0.880 ;
        RECT  1.490 0.460 1.590 1.775 ;
        RECT  1.590 0.570 1.610 1.775 ;
        RECT  1.610 1.635 2.260 1.775 ;
        RECT  1.610 0.570 2.260 0.730 ;
        RECT  11.810 0.470 12.070 0.590 ;
        RECT  11.690 0.470 11.810 1.550 ;
        RECT  10.760 0.470 11.690 0.590 ;
        RECT  11.610 1.060 11.690 1.280 ;
        RECT  10.600 0.470 10.760 1.570 ;
        RECT  12.230 1.910 12.470 2.070 ;
        RECT  10.350 1.910 12.230 2.050 ;
        RECT  10.210 0.620 10.350 2.050 ;
        RECT  10.190 0.620 10.210 1.740 ;
        RECT  12.950 1.060 13.090 1.280 ;
        RECT  12.830 1.060 12.950 1.790 ;
        RECT  11.090 1.670 12.830 1.790 ;
        RECT  11.090 0.710 11.190 0.850 ;
        RECT  10.970 0.710 11.090 1.790 ;
        RECT  10.130 1.520 10.190 1.740 ;
        RECT  10.470 1.410 10.600 1.570 ;
        RECT  10.910 1.370 10.970 1.590 ;
        RECT  11.280 1.420 11.310 1.540 ;
        RECT  8.620 1.050 8.700 1.270 ;
        RECT  9.380 1.410 9.570 1.810 ;
        RECT  7.990 0.470 8.140 1.730 ;
        RECT  5.330 1.400 5.420 1.560 ;
        RECT  7.620 1.470 7.710 1.690 ;
        RECT  4.530 1.550 4.640 1.710 ;
        RECT  4.920 1.410 5.050 1.570 ;
        RECT  5.710 1.400 5.830 1.540 ;
        RECT  3.070 1.050 3.150 1.270 ;
        RECT  3.830 1.410 3.970 1.810 ;
        RECT  2.400 0.470 2.520 1.650 ;
        RECT  0.550 1.595 0.770 2.015 ;
        RECT  1.350 1.615 1.490 1.775 ;
    END
END CMPE42D1

MACRO CMPE42D2
    CLASS CORE ;
    FOREIGN CMPE42D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.680 1.940 13.710 2.100 ;
        RECT  13.710 1.390 13.850 2.100 ;
        RECT  13.710 0.420 13.850 0.900 ;
        RECT  13.850 0.420 13.870 2.100 ;
        RECT  13.870 1.940 13.900 2.100 ;
        RECT  13.870 0.780 13.990 1.515 ;
        END
    END S
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 0.725 7.910 1.330 ;
        RECT  7.910 1.110 7.960 1.330 ;
        END
    END D
    PIN COX
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 1.410 7.130 1.550 ;
        RECT  6.980 0.450 7.130 0.870 ;
        RECT  7.130 0.450 7.200 1.550 ;
        RECT  7.200 0.750 7.270 1.550 ;
        END
    END COX
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.890 0.450 13.030 1.550 ;
        RECT  13.030 0.450 13.120 0.870 ;
        RECT  13.030 1.410 13.140 1.550 ;
        END
    END CO
    PIN CIX
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.050 1.080 12.250 1.235 ;
        RECT  12.250 1.005 12.710 1.235 ;
        END
    END CIX
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.180 1.035 6.490 1.195 ;
        RECT  6.490 1.005 6.950 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.970 1.830 1.515 ;
        RECT  1.830 0.970 1.860 1.210 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 14.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 14.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.300 1.670 6.795 1.790 ;
        RECT  6.795 1.670 6.915 2.050 ;
        RECT  6.915 1.930 7.550 2.050 ;
        RECT  7.550 1.930 7.770 2.100 ;
        RECT  7.770 1.930 8.460 2.050 ;
        RECT  8.460 0.710 8.600 2.050 ;
        RECT  8.600 1.400 8.630 2.050 ;
        RECT  8.600 0.710 8.710 0.850 ;
        RECT  7.605 1.650 7.920 1.810 ;
        RECT  7.605 0.450 7.920 0.605 ;
        RECT  4.380 0.620 4.400 1.710 ;
        RECT  4.400 0.620 4.540 2.050 ;
        RECT  4.540 1.910 6.420 2.050 ;
        RECT  6.420 1.910 6.660 2.070 ;
        RECT  4.790 0.470 4.950 1.570 ;
        RECT  5.800 1.060 5.910 1.280 ;
        RECT  4.950 0.470 5.910 0.590 ;
        RECT  5.910 0.470 6.050 1.550 ;
        RECT  6.050 0.470 6.260 0.590 ;
        RECT  6.260 0.450 6.480 0.870 ;
        RECT  6.050 1.410 6.490 1.550 ;
        RECT  5.500 0.760 5.620 1.540 ;
        RECT  5.620 1.420 5.710 1.540 ;
        RECT  5.620 0.760 5.790 0.900 ;
        RECT  2.890 1.050 2.910 2.050 ;
        RECT  2.910 0.760 3.030 2.050 ;
        RECT  3.030 0.760 3.150 0.920 ;
        RECT  3.030 1.930 3.960 2.050 ;
        RECT  3.960 1.530 4.030 2.050 ;
        RECT  3.990 0.620 4.030 0.860 ;
        RECT  4.030 0.620 4.080 2.050 ;
        RECT  4.080 0.620 4.150 1.750 ;
        RECT  3.650 0.450 3.710 0.950 ;
        RECT  3.710 0.450 3.790 1.810 ;
        RECT  3.790 0.450 3.830 1.550 ;
        RECT  3.830 1.040 3.910 1.260 ;
        RECT  2.260 0.470 2.360 0.660 ;
        RECT  2.260 1.490 2.380 1.650 ;
        RECT  2.360 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.530 1.275 ;
        RECT  3.530 1.055 3.590 1.275 ;
        RECT  0.420 0.460 0.640 0.880 ;
        RECT  0.640 1.895 0.810 2.015 ;
        RECT  0.640 0.760 0.810 0.880 ;
        RECT  0.810 0.760 0.930 2.015 ;
        RECT  0.930 1.060 1.060 1.280 ;
        RECT  0.930 1.895 2.540 2.015 ;
        RECT  2.540 0.710 2.680 2.015 ;
        RECT  2.680 1.470 2.710 2.015 ;
        RECT  2.680 0.710 2.780 0.850 ;
        RECT  1.110 0.460 1.230 0.880 ;
        RECT  1.230 0.460 1.330 1.775 ;
        RECT  1.330 0.570 1.350 1.775 ;
        RECT  1.350 1.635 2.000 1.775 ;
        RECT  1.350 0.570 2.000 0.730 ;
        RECT  5.300 0.710 5.380 0.850 ;
        RECT  5.180 0.710 5.300 1.790 ;
        RECT  5.160 0.710 5.180 0.850 ;
        RECT  9.380 1.045 9.540 1.275 ;
        RECT  9.330 1.045 9.380 1.165 ;
        RECT  9.210 0.470 9.330 1.165 ;
        RECT  8.280 0.470 9.210 0.590 ;
        RECT  8.150 0.470 8.280 1.710 ;
        RECT  8.120 0.470 8.150 0.750 ;
        RECT  9.800 1.040 9.880 1.260 ;
        RECT  9.710 0.470 9.800 1.550 ;
        RECT  9.680 0.470 9.710 1.810 ;
        RECT  9.550 0.470 9.680 0.690 ;
        RECT  10.000 0.640 10.120 1.880 ;
        RECT  9.930 0.640 10.000 0.860 ;
        RECT  9.880 1.660 10.000 2.050 ;
        RECT  8.950 1.930 9.880 2.050 ;
        RECT  8.950 0.710 9.070 0.870 ;
        RECT  8.830 0.710 8.950 2.050 ;
        RECT  8.810 1.050 8.830 2.050 ;
        RECT  11.540 0.730 11.660 0.950 ;
        RECT  11.540 1.420 11.630 1.540 ;
        RECT  11.420 0.730 11.540 1.540 ;
        RECT  11.920 1.410 12.410 1.550 ;
        RECT  12.180 0.450 12.400 0.870 ;
        RECT  11.920 0.470 12.180 0.590 ;
        RECT  11.800 0.470 11.920 1.550 ;
        RECT  10.870 0.470 11.800 0.590 ;
        RECT  11.720 1.060 11.800 1.280 ;
        RECT  10.710 0.470 10.870 1.570 ;
        RECT  12.340 1.910 12.580 2.070 ;
        RECT  10.460 1.910 12.340 2.050 ;
        RECT  10.320 0.620 10.460 2.050 ;
        RECT  10.300 0.620 10.320 1.740 ;
        RECT  13.430 1.080 13.720 1.240 ;
        RECT  13.310 1.080 13.430 1.790 ;
        RECT  11.200 1.670 13.310 1.790 ;
        RECT  11.200 0.710 11.300 0.850 ;
        RECT  11.080 0.710 11.200 1.790 ;
        RECT  11.020 1.370 11.080 1.590 ;
        RECT  10.240 1.520 10.300 1.740 ;
        RECT  10.580 1.410 10.710 1.570 ;
        RECT  11.390 1.420 11.420 1.540 ;
        RECT  8.730 1.050 8.810 1.270 ;
        RECT  9.490 1.410 9.680 1.810 ;
        RECT  8.090 1.490 8.150 1.710 ;
        RECT  5.070 1.400 5.180 1.560 ;
        RECT  7.485 0.450 7.605 1.810 ;
        RECT  4.270 1.550 4.380 1.710 ;
        RECT  4.660 1.410 4.790 1.570 ;
        RECT  5.470 1.420 5.500 1.540 ;
        RECT  2.810 1.050 2.890 1.270 ;
        RECT  3.570 1.410 3.710 1.810 ;
        RECT  2.140 0.470 2.260 1.650 ;
        RECT  0.420 1.615 0.640 2.015 ;
        RECT  1.090 1.615 1.230 1.775 ;
    END
END CMPE42D2

MACRO DCAP
    CLASS CORE ;
    FOREIGN DCAP 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.360 0.420 0.580 0.830 ;
        RECT  0.080 0.670 0.240 1.440 ;
        RECT  0.400 0.950 0.560 2.090 ;
        RECT  0.240 0.670 0.360 0.830 ;
    END
END DCAP

MACRO DCAP16
    CLASS CORE ;
    FOREIGN DCAP16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.840 0.420 5.060 0.830 ;
        RECT  4.730 0.710 4.840 0.830 ;
        RECT  4.230 1.240 4.610 1.400 ;
        RECT  4.870 0.950 5.040 2.090 ;
        RECT  4.610 0.710 4.730 1.400 ;
    END
END DCAP16

MACRO DCAP32
    CLASS CORE ;
    FOREIGN DCAP32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.960 0.420 10.180 0.830 ;
        RECT  9.850 0.710 9.960 0.830 ;
        RECT  9.350 1.240 9.730 1.400 ;
        RECT  9.990 0.950 10.160 2.090 ;
        RECT  9.730 0.710 9.850 1.400 ;
    END
END DCAP32

MACRO DCAP4
    CLASS CORE ;
    FOREIGN DCAP4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.000 0.420 1.220 0.830 ;
        RECT  0.890 0.710 1.000 0.830 ;
        RECT  0.390 1.240 0.770 1.400 ;
        RECT  1.030 0.950 1.200 2.090 ;
        RECT  0.770 0.710 0.890 1.400 ;
    END
END DCAP4

MACRO DCAP64
    CLASS CORE ;
    FOREIGN DCAP64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 20.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 20.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  20.200 0.420 20.420 0.830 ;
        RECT  20.090 0.710 20.200 0.830 ;
        RECT  19.590 1.240 19.970 1.400 ;
        RECT  20.230 0.950 20.400 2.090 ;
        RECT  19.970 0.710 20.090 1.400 ;
    END
END DCAP64

MACRO DCAP8
    CLASS CORE ;
    FOREIGN DCAP8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 0.420 2.500 0.830 ;
        RECT  2.170 0.710 2.280 0.830 ;
        RECT  1.670 1.240 2.050 1.400 ;
        RECT  2.310 0.950 2.480 2.090 ;
        RECT  2.050 0.710 2.170 1.400 ;
    END
END DCAP8

MACRO DEL0
    CLASS CORE ;
    FOREIGN DEL0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.660 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.820 0.730 0.980 1.760 ;
        RECT  0.280 0.730 0.820 0.850 ;
        RECT  0.280 1.640 0.820 1.760 ;
        RECT  0.060 0.430 0.280 0.850 ;
        RECT  1.350 1.080 2.100 1.240 ;
        RECT  1.350 1.960 1.380 2.100 ;
        RECT  1.190 0.420 1.350 2.100 ;
        RECT  2.470 1.050 2.510 1.270 ;
        RECT  2.350 0.780 2.470 1.510 ;
        RECT  1.690 0.780 2.350 0.900 ;
        RECT  1.690 1.390 2.350 1.510 ;
        RECT  1.690 1.960 1.720 2.100 ;
        RECT  1.530 0.420 1.690 0.900 ;
        RECT  1.530 1.390 1.690 2.100 ;
        RECT  1.500 1.960 1.530 2.100 ;
        RECT  1.160 1.960 1.190 2.100 ;
        RECT  0.060 1.640 0.280 2.060 ;
    END
END DEL0

MACRO DEL01
    CLASS CORE ;
    FOREIGN DEL01 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.940 2.630 2.100 ;
        RECT  2.630 1.390 2.650 2.100 ;
        RECT  2.650 0.440 2.790 2.100 ;
        RECT  2.790 1.940 2.820 2.100 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.765 0.700 1.775 ;
        RECT  0.280 0.765 0.560 0.885 ;
        RECT  0.280 1.655 0.560 1.775 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  1.340 1.050 1.410 1.270 ;
        RECT  2.390 0.470 2.530 1.290 ;
        RECT  1.680 0.470 2.390 0.590 ;
        RECT  1.900 0.720 2.060 1.890 ;
        RECT  1.180 0.440 1.340 1.890 ;
        RECT  0.820 0.440 0.960 1.890 ;
        RECT  0.060 1.655 0.280 2.075 ;
        RECT  1.530 0.460 1.680 1.890 ;
    END
END DEL01

MACRO DEL015
    CLASS CORE ;
    FOREIGN DEL015 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.940 3.210 2.100 ;
        RECT  3.210 1.390 3.290 2.100 ;
        RECT  3.210 0.440 3.290 0.940 ;
        RECT  3.290 0.440 3.370 2.100 ;
        RECT  3.370 1.940 3.400 2.100 ;
        RECT  3.370 0.820 3.430 1.515 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.780 0.300 ;
        RECT  2.780 -0.300 3.000 0.340 ;
        RECT  3.000 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.780 2.820 ;
        RECT  2.780 2.180 3.000 2.820 ;
        RECT  3.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.630 0.765 0.790 1.775 ;
        RECT  0.280 0.765 0.630 0.885 ;
        RECT  0.280 1.655 0.630 1.775 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  1.570 1.050 1.660 1.270 ;
        RECT  2.880 0.470 3.040 1.290 ;
        RECT  1.940 0.470 2.880 0.590 ;
        RECT  2.160 0.710 2.320 1.890 ;
        RECT  1.410 0.435 1.570 1.890 ;
        RECT  1.030 0.435 1.190 1.890 ;
        RECT  0.060 1.655 0.280 2.075 ;
        RECT  1.780 0.470 1.940 1.890 ;
    END
END DEL015

MACRO DEL02
    CLASS CORE ;
    FOREIGN DEL02 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.940 3.210 2.100 ;
        RECT  3.210 1.390 3.290 2.100 ;
        RECT  3.210 0.440 3.290 0.940 ;
        RECT  3.290 0.440 3.370 2.100 ;
        RECT  3.370 1.940 3.400 2.100 ;
        RECT  3.370 0.820 3.430 1.515 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 2.780 0.300 ;
        RECT  2.780 -0.300 3.000 0.340 ;
        RECT  3.000 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 2.780 2.820 ;
        RECT  2.780 2.180 3.000 2.820 ;
        RECT  3.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.630 0.765 0.790 1.775 ;
        RECT  0.280 0.765 0.630 0.885 ;
        RECT  0.280 1.655 0.630 1.775 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  1.570 1.050 1.660 1.270 ;
        RECT  2.880 0.470 3.040 1.290 ;
        RECT  1.940 0.470 2.880 0.590 ;
        RECT  2.160 0.710 2.320 1.630 ;
        RECT  1.410 0.675 1.570 1.630 ;
        RECT  1.030 0.675 1.190 1.630 ;
        RECT  0.060 1.655 0.280 2.075 ;
        RECT  1.780 0.470 1.940 1.630 ;
    END
END DEL02

MACRO DEL1
    CLASS CORE ;
    FOREIGN DEL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.960 3.270 2.100 ;
        RECT  3.270 0.660 3.430 2.100 ;
        RECT  3.430 1.960 3.460 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 1.080 1.330 1.240 ;
        RECT  0.830 0.730 0.950 1.760 ;
        RECT  0.280 0.730 0.830 0.850 ;
        RECT  0.280 1.640 0.830 1.760 ;
        RECT  0.060 0.430 0.280 0.850 ;
        RECT  1.670 1.080 2.700 1.240 ;
        RECT  1.670 1.960 1.700 2.100 ;
        RECT  1.510 0.660 1.670 2.100 ;
        RECT  3.130 1.040 3.150 1.260 ;
        RECT  2.990 0.710 3.130 1.510 ;
        RECT  1.800 0.710 2.990 0.870 ;
        RECT  2.010 1.390 2.990 1.510 ;
        RECT  2.010 1.960 2.040 2.100 ;
        RECT  1.850 1.390 2.010 2.100 ;
        RECT  1.820 1.960 1.850 2.100 ;
        RECT  1.480 1.960 1.510 2.100 ;
        RECT  0.060 1.640 0.280 2.060 ;
    END
END DEL1

MACRO DEL2
    CLASS CORE ;
    FOREIGN DEL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.960 4.230 2.100 ;
        RECT  4.230 0.670 4.390 2.100 ;
        RECT  4.390 1.960 4.420 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.060 1.080 1.700 1.240 ;
        RECT  0.940 0.730 1.060 1.760 ;
        RECT  0.280 0.730 0.940 0.850 ;
        RECT  0.280 1.640 0.940 1.760 ;
        RECT  0.060 0.430 0.280 0.850 ;
        RECT  2.150 1.080 3.560 1.240 ;
        RECT  2.150 1.960 2.180 2.100 ;
        RECT  1.990 0.620 2.150 2.100 ;
        RECT  3.950 0.810 4.110 1.510 ;
        RECT  2.490 0.810 3.950 0.930 ;
        RECT  2.490 1.390 3.950 1.510 ;
        RECT  2.490 1.960 2.520 2.100 ;
        RECT  2.330 0.430 2.490 0.930 ;
        RECT  2.330 1.390 2.490 2.100 ;
        RECT  2.300 1.960 2.330 2.100 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  0.060 1.640 0.280 2.060 ;
    END
END DEL2

MACRO DEL3
    CLASS CORE ;
    FOREIGN DEL3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.840 1.960 4.870 2.100 ;
        RECT  4.870 0.670 5.030 2.100 ;
        RECT  5.030 1.960 5.060 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.085 1.080 1.985 1.240 ;
        RECT  0.965 0.730 1.085 1.760 ;
        RECT  0.280 0.730 0.965 0.850 ;
        RECT  0.280 1.640 0.965 1.760 ;
        RECT  0.060 0.430 0.280 0.850 ;
        RECT  2.470 1.080 4.175 1.240 ;
        RECT  2.470 1.960 2.500 2.100 ;
        RECT  2.310 0.620 2.470 2.100 ;
        RECT  4.710 1.050 4.750 1.270 ;
        RECT  4.590 0.780 4.710 1.510 ;
        RECT  2.810 0.780 4.590 0.900 ;
        RECT  2.810 1.390 4.590 1.510 ;
        RECT  2.810 1.960 2.840 2.100 ;
        RECT  2.650 0.420 2.810 0.900 ;
        RECT  2.650 1.390 2.810 2.100 ;
        RECT  2.620 1.960 2.650 2.100 ;
        RECT  2.280 1.960 2.310 2.100 ;
        RECT  0.060 1.640 0.280 2.060 ;
    END
END DEL3

MACRO DEL4
    CLASS CORE ;
    FOREIGN DEL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 1.960 5.510 2.100 ;
        RECT  5.510 0.670 5.670 2.100 ;
        RECT  5.670 1.960 5.700 2.100 ;
        END
    END Z
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 5.080 0.300 ;
        RECT  5.080 -0.300 5.300 0.340 ;
        RECT  5.300 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.130 1.080 2.290 1.240 ;
        RECT  1.010 0.760 1.130 1.760 ;
        RECT  0.290 0.760 1.010 0.880 ;
        RECT  0.290 1.640 1.010 1.760 ;
        RECT  0.070 0.430 0.290 0.880 ;
        RECT  2.790 1.080 4.770 1.240 ;
        RECT  2.790 1.960 2.820 2.100 ;
        RECT  2.630 0.630 2.790 2.100 ;
        RECT  5.230 0.780 5.390 1.510 ;
        RECT  3.130 0.780 5.230 0.900 ;
        RECT  3.130 1.390 5.230 1.510 ;
        RECT  3.130 1.960 3.160 2.100 ;
        RECT  2.970 0.420 3.130 0.900 ;
        RECT  2.970 1.390 3.130 2.100 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  0.070 1.640 0.290 2.060 ;
        RECT  2.940 1.960 2.970 2.100 ;
    END
END DEL4

MACRO DFCND1
    CLASS CORE ;
    FOREIGN DFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.940 6.790 2.100 ;
        RECT  6.790 0.420 6.950 2.100 ;
        RECT  6.950 1.940 6.980 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.920 1.940 5.950 2.100 ;
        RECT  5.950 1.390 6.110 2.100 ;
        RECT  6.110 1.940 6.140 2.100 ;
        RECT  6.110 1.390 6.170 1.515 ;
        RECT  5.900 0.710 6.170 0.830 ;
        RECT  6.170 0.710 6.310 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.710 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.285 4.970 1.515 ;
        RECT  4.970 1.190 5.130 1.515 ;
        RECT  5.130 1.285 5.350 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.000 0.300 ;
        RECT  1.000 -0.300 1.220 0.480 ;
        RECT  1.220 -0.300 2.720 0.300 ;
        RECT  2.720 -0.300 2.880 0.720 ;
        RECT  2.880 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.550 ;
        RECT  5.000 -0.300 6.340 0.300 ;
        RECT  6.340 -0.300 6.560 0.340 ;
        RECT  6.560 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.040 2.820 ;
        RECT  1.040 2.030 1.260 2.820 ;
        RECT  1.260 2.220 2.480 2.820 ;
        RECT  2.480 2.030 2.700 2.820 ;
        RECT  2.700 2.220 3.110 2.820 ;
        RECT  3.110 1.670 3.330 2.820 ;
        RECT  3.330 2.220 4.670 2.820 ;
        RECT  4.670 2.180 4.890 2.820 ;
        RECT  4.890 2.220 5.500 2.820 ;
        RECT  5.500 2.180 5.720 2.820 ;
        RECT  5.720 2.220 6.340 2.820 ;
        RECT  6.340 2.180 6.560 2.820 ;
        RECT  6.560 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.900 1.120 4.060 2.050 ;
        RECT  4.060 1.930 5.530 2.050 ;
        RECT  5.530 1.190 5.690 2.050 ;
        RECT  0.730 0.710 0.960 0.870 ;
        RECT  0.960 0.710 1.120 1.730 ;
        RECT  1.120 0.710 1.390 0.830 ;
        RECT  1.390 0.470 1.530 0.830 ;
        RECT  1.530 0.470 2.290 0.590 ;
        RECT  2.290 0.470 2.410 0.960 ;
        RECT  2.410 0.840 3.000 0.960 ;
        RECT  3.000 0.470 3.120 0.960 ;
        RECT  3.120 0.470 4.080 0.590 ;
        RECT  4.080 0.430 4.300 0.590 ;
        RECT  3.240 0.710 3.340 0.930 ;
        RECT  3.340 0.710 3.460 1.540 ;
        RECT  3.460 1.420 3.520 1.540 ;
        RECT  3.520 1.420 3.680 1.840 ;
        RECT  1.690 0.740 1.830 0.900 ;
        RECT  1.830 0.740 1.950 1.830 ;
        RECT  1.950 1.080 3.220 1.200 ;
        RECT  0.060 0.705 0.420 0.865 ;
        RECT  0.420 0.705 0.540 2.050 ;
        RECT  0.540 1.910 0.620 2.050 ;
        RECT  0.620 1.910 0.860 2.070 ;
        RECT  3.780 1.120 3.900 1.240 ;
        RECT  5.890 0.950 6.050 1.270 ;
        RECT  5.610 0.950 5.890 1.070 ;
        RECT  5.450 0.710 5.610 1.070 ;
        RECT  4.770 0.950 5.450 1.070 ;
        RECT  4.770 1.650 5.330 1.810 ;
        RECT  6.510 0.470 6.670 1.290 ;
        RECT  5.300 0.470 6.510 0.590 ;
        RECT  5.180 0.470 5.300 0.830 ;
        RECT  4.510 0.670 5.180 0.830 ;
        RECT  4.390 0.670 4.510 1.810 ;
        RECT  3.950 0.830 4.390 0.990 ;
        RECT  4.240 1.650 4.390 1.810 ;
        RECT  4.630 0.950 4.770 1.810 ;
        RECT  3.620 0.770 3.780 1.240 ;
        RECT  0.730 1.570 0.960 1.730 ;
        RECT  2.280 1.380 3.340 1.540 ;
        RECT  1.680 1.670 1.830 1.830 ;
        RECT  2.080 1.670 2.970 1.830 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFCND1

MACRO DFCND2
    CLASS CORE ;
    FOREIGN DFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.250 1.940 7.280 2.100 ;
        RECT  7.280 1.390 7.440 2.100 ;
        RECT  7.280 0.420 7.440 0.900 ;
        RECT  7.440 1.390 7.450 1.515 ;
        RECT  7.440 0.780 7.450 0.900 ;
        RECT  7.440 1.940 7.470 2.100 ;
        RECT  7.450 0.780 7.590 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.420 1.940 6.450 2.100 ;
        RECT  6.450 1.390 6.490 2.100 ;
        RECT  6.400 0.740 6.490 0.900 ;
        RECT  6.490 0.740 6.610 2.100 ;
        RECT  6.610 1.940 6.640 2.100 ;
        RECT  6.610 0.740 6.640 1.530 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.020 1.700 1.240 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.285 4.920 1.515 ;
        RECT  4.920 1.190 5.080 1.515 ;
        RECT  5.080 1.285 5.350 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.020 0.300 ;
        RECT  1.020 -0.300 1.240 0.480 ;
        RECT  1.240 -0.300 2.690 0.300 ;
        RECT  2.690 -0.300 2.830 0.740 ;
        RECT  2.830 -0.300 4.730 0.300 ;
        RECT  4.730 -0.300 4.950 0.550 ;
        RECT  4.950 -0.300 6.020 0.300 ;
        RECT  6.020 -0.300 6.240 0.340 ;
        RECT  6.240 -0.300 6.840 0.300 ;
        RECT  6.840 -0.300 7.060 0.340 ;
        RECT  7.060 -0.300 7.650 0.300 ;
        RECT  7.650 -0.300 7.870 0.340 ;
        RECT  7.870 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.010 2.820 ;
        RECT  1.010 2.030 1.230 2.820 ;
        RECT  1.230 2.220 2.430 2.820 ;
        RECT  2.430 2.030 2.650 2.820 ;
        RECT  2.650 2.220 3.060 2.820 ;
        RECT  3.060 1.670 3.280 2.820 ;
        RECT  3.280 2.220 4.620 2.820 ;
        RECT  4.620 2.180 4.840 2.820 ;
        RECT  4.840 2.220 6.840 2.820 ;
        RECT  6.840 2.180 7.060 2.820 ;
        RECT  7.060 2.220 7.650 2.820 ;
        RECT  7.650 2.180 7.870 2.820 ;
        RECT  7.870 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.470 1.420 3.630 1.970 ;
        RECT  1.790 1.410 1.830 1.835 ;
        RECT  1.710 0.730 1.830 0.890 ;
        RECT  1.830 0.730 1.910 1.835 ;
        RECT  1.910 0.730 1.950 1.545 ;
        RECT  1.950 1.100 3.170 1.240 ;
        RECT  0.060 0.445 0.420 0.605 ;
        RECT  0.420 0.445 0.540 1.750 ;
        RECT  0.540 1.055 0.730 1.275 ;
        RECT  3.410 1.420 3.470 1.540 ;
        RECT  3.290 0.710 3.410 1.540 ;
        RECT  3.190 0.710 3.290 0.930 ;
        RECT  4.030 0.430 4.250 0.590 ;
        RECT  3.070 0.470 4.030 0.590 ;
        RECT  2.950 0.470 3.070 0.980 ;
        RECT  2.220 0.860 2.950 0.980 ;
        RECT  2.100 0.470 2.220 0.980 ;
        RECT  1.520 0.470 2.100 0.590 ;
        RECT  1.400 0.470 1.520 0.830 ;
        RECT  1.120 0.710 1.400 0.830 ;
        RECT  0.965 0.710 1.120 1.635 ;
        RECT  0.730 0.710 0.965 0.870 ;
        RECT  5.480 1.190 5.640 2.050 ;
        RECT  4.010 1.930 5.480 2.050 ;
        RECT  3.850 1.120 4.010 2.050 ;
        RECT  3.730 1.120 3.850 1.240 ;
        RECT  5.920 1.050 6.370 1.270 ;
        RECT  5.760 0.950 5.920 1.960 ;
        RECT  5.560 0.950 5.760 1.070 ;
        RECT  5.400 0.710 5.560 1.070 ;
        RECT  4.740 0.950 5.400 1.070 ;
        RECT  4.740 1.650 5.270 1.810 ;
        RECT  7.030 1.080 7.320 1.240 ;
        RECT  6.890 0.470 7.030 1.240 ;
        RECT  5.250 0.470 6.890 0.590 ;
        RECT  5.130 0.470 5.250 0.830 ;
        RECT  4.460 0.670 5.130 0.830 ;
        RECT  4.340 0.670 4.460 1.810 ;
        RECT  3.900 0.810 4.340 0.970 ;
        RECT  4.580 0.950 4.740 1.810 ;
        RECT  4.190 1.650 4.340 1.810 ;
        RECT  3.570 0.760 3.730 1.240 ;
        RECT  0.730 1.475 0.965 1.635 ;
        RECT  2.230 1.380 3.290 1.540 ;
        RECT  1.630 1.675 1.790 1.835 ;
        RECT  2.030 1.670 2.920 1.830 ;
        RECT  0.060 1.590 0.420 1.750 ;
    END
END DFCND2

MACRO DFCND4
    CLASS CORE ;
    FOREIGN DFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.590 1.650 8.910 2.030 ;
        RECT  8.590 0.490 8.910 0.870 ;
        RECT  8.910 0.490 9.330 2.030 ;
        RECT  9.330 1.650 9.500 2.030 ;
        RECT  9.330 0.490 9.500 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 1.650 7.310 2.030 ;
        RECT  7.210 0.760 7.310 0.920 ;
        RECT  7.310 0.760 7.730 2.030 ;
        RECT  7.730 1.650 8.120 2.030 ;
        RECT  7.730 0.760 8.140 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.830 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.050 1.190 6.210 1.515 ;
        RECT  6.210 1.285 6.630 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.480 ;
        RECT  1.370 -0.300 2.810 0.300 ;
        RECT  2.810 -0.300 2.970 0.720 ;
        RECT  2.970 -0.300 4.880 0.300 ;
        RECT  4.880 -0.300 5.100 0.550 ;
        RECT  5.100 -0.300 6.180 0.300 ;
        RECT  6.180 -0.300 6.400 0.340 ;
        RECT  6.400 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.060 2.820 ;
        RECT  1.060 2.000 1.280 2.820 ;
        RECT  1.280 2.220 2.570 2.820 ;
        RECT  2.570 2.030 2.790 2.820 ;
        RECT  2.790 2.220 3.200 2.820 ;
        RECT  3.200 1.670 3.420 2.820 ;
        RECT  3.420 2.220 4.760 2.820 ;
        RECT  4.760 2.180 4.980 2.820 ;
        RECT  4.980 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.105 0.790 1.265 ;
        RECT  0.420 0.725 0.540 1.795 ;
        RECT  0.280 0.725 0.420 0.885 ;
        RECT  0.280 1.635 0.420 1.795 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  2.080 1.080 3.310 1.240 ;
        RECT  2.010 0.710 2.080 1.505 ;
        RECT  1.960 0.710 2.010 1.830 ;
        RECT  1.910 0.710 1.960 0.930 ;
        RECT  1.890 1.385 1.960 1.830 ;
        RECT  3.610 1.420 3.770 1.970 ;
        RECT  3.550 1.420 3.610 1.540 ;
        RECT  3.430 0.710 3.550 1.540 ;
        RECT  3.330 0.710 3.430 0.930 ;
        RECT  4.170 0.430 4.390 0.590 ;
        RECT  3.210 0.470 4.170 0.590 ;
        RECT  3.090 0.470 3.210 0.960 ;
        RECT  2.515 0.840 3.090 0.960 ;
        RECT  2.395 0.470 2.515 0.960 ;
        RECT  1.710 0.470 2.395 0.590 ;
        RECT  1.570 0.470 1.710 0.720 ;
        RECT  1.240 0.600 1.570 0.720 ;
        RECT  1.090 0.600 1.240 1.695 ;
        RECT  0.780 0.600 1.090 0.760 ;
        RECT  5.510 1.190 5.660 2.050 ;
        RECT  5.500 1.190 5.510 1.410 ;
        RECT  4.150 1.930 5.510 2.050 ;
        RECT  3.990 1.120 4.150 2.050 ;
        RECT  3.870 1.120 3.990 1.240 ;
        RECT  6.630 0.950 6.850 1.160 ;
        RECT  5.930 0.950 6.630 1.070 ;
        RECT  5.930 1.685 6.090 2.100 ;
        RECT  5.870 0.950 5.930 2.100 ;
        RECT  5.780 0.950 5.870 1.845 ;
        RECT  5.720 0.950 5.780 1.070 ;
        RECT  5.560 0.710 5.720 1.070 ;
        RECT  4.880 0.950 5.560 1.070 ;
        RECT  4.880 1.650 5.390 1.810 ;
        RECT  8.400 1.080 8.690 1.240 ;
        RECT  8.280 0.470 8.400 1.240 ;
        RECT  7.090 0.470 8.280 0.590 ;
        RECT  6.970 0.470 7.090 1.845 ;
        RECT  6.740 0.470 6.970 0.590 ;
        RECT  6.740 1.685 6.970 1.845 ;
        RECT  6.520 0.470 6.740 0.650 ;
        RECT  6.520 1.685 6.740 2.100 ;
        RECT  5.410 0.470 6.520 0.590 ;
        RECT  5.290 0.470 5.410 0.830 ;
        RECT  4.600 0.670 5.290 0.830 ;
        RECT  4.480 0.670 4.600 1.810 ;
        RECT  4.040 0.810 4.480 0.970 ;
        RECT  4.720 0.950 4.880 1.810 ;
        RECT  3.710 0.760 3.870 1.240 ;
        RECT  4.330 1.650 4.480 1.810 ;
        RECT  0.780 1.535 1.090 1.695 ;
        RECT  2.370 1.380 3.430 1.540 ;
        RECT  1.770 1.670 1.890 1.830 ;
        RECT  2.150 1.670 3.060 1.830 ;
        RECT  0.060 1.635 0.280 2.055 ;
        LAYER M1 ;
        RECT  8.590 1.650 8.695 2.030 ;
        RECT  8.590 0.490 8.695 0.870 ;
        RECT  7.945 1.650 8.120 2.030 ;
        RECT  7.945 0.760 8.140 0.920 ;
    END
END DFCND4

MACRO DFCNQD1
    CLASS CORE ;
    FOREIGN DFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.720 1.940 5.750 2.100 ;
        RECT  5.750 1.390 5.910 2.100 ;
        RECT  5.910 1.940 5.940 2.100 ;
        RECT  5.720 0.420 5.940 0.830 ;
        RECT  5.910 1.390 6.170 1.515 ;
        RECT  5.940 0.710 6.170 0.830 ;
        RECT  6.170 0.710 6.310 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.680 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.285 4.910 1.515 ;
        RECT  4.910 1.190 5.070 1.515 ;
        RECT  5.070 1.285 5.350 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.000 0.300 ;
        RECT  1.000 -0.300 1.220 0.480 ;
        RECT  1.220 -0.300 2.660 0.300 ;
        RECT  2.660 -0.300 2.820 0.520 ;
        RECT  2.820 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.940 0.830 ;
        RECT  4.940 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.000 2.820 ;
        RECT  1.000 2.000 1.220 2.820 ;
        RECT  1.220 2.220 2.420 2.820 ;
        RECT  2.420 2.030 2.640 2.820 ;
        RECT  2.640 2.220 3.050 2.820 ;
        RECT  3.050 1.670 3.270 2.820 ;
        RECT  3.270 2.220 4.610 2.820 ;
        RECT  4.610 2.180 4.830 2.820 ;
        RECT  4.830 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.190 0.640 2.940 0.760 ;
        RECT  2.940 0.470 3.060 0.760 ;
        RECT  3.060 0.470 4.020 0.590 ;
        RECT  4.020 0.430 4.240 0.590 ;
        RECT  3.180 0.710 3.340 1.505 ;
        RECT  3.340 1.385 3.460 1.505 ;
        RECT  3.460 1.385 3.620 1.840 ;
        RECT  1.760 0.710 1.800 0.930 ;
        RECT  1.800 0.710 1.830 1.820 ;
        RECT  1.830 0.710 1.920 1.550 ;
        RECT  1.920 1.000 1.930 1.550 ;
        RECT  1.930 1.000 3.060 1.160 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 2.050 ;
        RECT  0.540 1.910 0.620 2.050 ;
        RECT  0.620 1.910 0.860 2.070 ;
        RECT  2.070 0.470 2.190 0.760 ;
        RECT  1.540 0.470 2.070 0.590 ;
        RECT  1.420 0.470 1.540 0.800 ;
        RECT  0.940 0.680 1.420 0.800 ;
        RECT  0.940 1.080 1.120 1.300 ;
        RECT  4.450 0.670 4.570 0.830 ;
        RECT  4.330 0.670 4.450 1.810 ;
        RECT  3.890 0.830 4.330 0.990 ;
        RECT  5.490 1.190 5.630 1.770 ;
        RECT  5.470 1.190 5.490 2.050 ;
        RECT  5.370 1.650 5.470 2.050 ;
        RECT  4.000 1.930 5.370 2.050 ;
        RECT  3.840 1.120 4.000 2.050 ;
        RECT  3.720 1.120 3.840 1.240 ;
        RECT  5.890 0.950 6.050 1.270 ;
        RECT  5.550 0.950 5.890 1.070 ;
        RECT  5.390 0.650 5.550 1.070 ;
        RECT  4.730 0.950 5.390 1.070 ;
        RECT  4.730 1.650 5.250 1.810 ;
        RECT  4.570 0.950 4.730 1.810 ;
        RECT  3.560 0.770 3.720 1.240 ;
        RECT  4.180 1.650 4.330 1.810 ;
        RECT  0.780 0.680 0.940 1.780 ;
        RECT  2.220 1.345 3.180 1.505 ;
        RECT  1.670 1.430 1.800 1.820 ;
        RECT  2.000 1.650 2.910 1.815 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFCNQD1

MACRO DFCNQD2
    CLASS CORE ;
    FOREIGN DFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.600 6.570 2.020 ;
        RECT  6.350 0.490 6.570 0.910 ;
        RECT  6.570 1.600 6.810 1.760 ;
        RECT  6.570 0.725 6.810 0.910 ;
        RECT  6.810 0.725 6.950 1.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.680 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.990 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.005 5.990 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.010 0.300 ;
        RECT  1.010 -0.300 1.230 0.490 ;
        RECT  1.230 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.830 0.740 ;
        RECT  2.830 -0.300 4.670 0.300 ;
        RECT  4.670 -0.300 4.890 0.490 ;
        RECT  4.890 -0.300 5.955 0.300 ;
        RECT  5.955 -0.300 6.175 0.340 ;
        RECT  6.175 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.010 2.820 ;
        RECT  1.010 2.000 1.230 2.820 ;
        RECT  1.230 2.220 2.430 2.820 ;
        RECT  2.430 2.030 2.650 2.820 ;
        RECT  2.650 2.220 3.060 2.820 ;
        RECT  3.060 1.670 3.280 2.820 ;
        RECT  3.280 2.220 4.515 2.820 ;
        RECT  4.515 2.180 4.735 2.820 ;
        RECT  4.735 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.020 0.770 1.180 ;
        RECT  0.420 0.705 0.540 1.850 ;
        RECT  0.060 0.705 0.420 0.865 ;
        RECT  1.950 1.100 3.170 1.260 ;
        RECT  1.930 0.760 1.950 1.260 ;
        RECT  1.900 0.760 1.930 1.535 ;
        RECT  1.810 0.760 1.900 1.830 ;
        RECT  1.710 0.760 1.810 0.920 ;
        RECT  1.780 1.385 1.810 1.830 ;
        RECT  3.470 1.420 3.630 1.970 ;
        RECT  3.410 1.420 3.470 1.540 ;
        RECT  3.290 0.710 3.410 1.540 ;
        RECT  3.190 0.710 3.290 0.930 ;
        RECT  4.010 0.430 4.250 0.590 ;
        RECT  3.070 0.470 4.010 0.590 ;
        RECT  2.950 0.470 3.070 0.980 ;
        RECT  2.480 0.860 2.950 0.980 ;
        RECT  2.360 0.470 2.480 0.980 ;
        RECT  1.490 0.470 2.360 0.590 ;
        RECT  1.370 0.470 1.490 0.830 ;
        RECT  1.110 0.710 1.370 0.830 ;
        RECT  0.950 0.710 1.110 1.570 ;
        RECT  0.730 0.710 0.950 0.870 ;
        RECT  5.310 1.190 5.470 2.050 ;
        RECT  4.010 1.930 5.310 2.050 ;
        RECT  3.850 1.120 4.010 2.050 ;
        RECT  3.730 1.120 3.850 1.240 ;
        RECT  6.230 1.080 6.460 1.240 ;
        RECT  6.110 0.720 6.230 1.240 ;
        RECT  5.710 0.720 6.110 0.840 ;
        RECT  5.710 1.780 5.900 1.940 ;
        RECT  5.590 0.720 5.710 1.940 ;
        RECT  5.500 0.720 5.590 1.070 ;
        RECT  5.340 0.680 5.500 1.070 ;
        RECT  5.130 0.950 5.340 1.070 ;
        RECT  5.130 1.650 5.190 1.810 ;
        RECT  4.970 0.950 5.130 1.810 ;
        RECT  3.570 0.760 3.730 1.240 ;
        RECT  3.900 0.810 4.590 0.970 ;
        RECT  0.730 1.410 0.950 1.570 ;
        RECT  2.230 1.380 3.290 1.540 ;
        RECT  1.630 1.670 1.780 1.830 ;
        RECT  2.030 1.670 2.920 1.830 ;
        RECT  0.060 1.690 0.420 1.850 ;
        RECT  4.480 1.220 4.970 1.380 ;
    END
END DFCNQD2

MACRO DFCNQD4
    CLASS CORE ;
    FOREIGN DFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.650 6.670 2.030 ;
        RECT  6.350 0.490 6.670 0.870 ;
        RECT  6.670 0.490 7.090 2.030 ;
        RECT  7.090 1.650 7.260 2.030 ;
        RECT  7.090 0.490 7.260 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.690 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.990 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.830 1.005 5.990 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.020 0.300 ;
        RECT  1.020 -0.300 1.240 0.490 ;
        RECT  1.240 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.830 0.740 ;
        RECT  2.830 -0.300 4.670 0.300 ;
        RECT  4.670 -0.300 4.890 0.520 ;
        RECT  4.890 -0.300 5.955 0.300 ;
        RECT  5.955 -0.300 6.175 0.340 ;
        RECT  6.175 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.010 2.820 ;
        RECT  1.010 2.000 1.230 2.820 ;
        RECT  1.230 2.220 2.430 2.820 ;
        RECT  2.430 2.030 2.650 2.820 ;
        RECT  2.650 2.220 3.060 2.820 ;
        RECT  3.060 1.670 3.280 2.820 ;
        RECT  3.280 2.220 4.515 2.820 ;
        RECT  4.515 2.180 4.735 2.820 ;
        RECT  4.735 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.020 0.770 1.180 ;
        RECT  0.420 0.660 0.540 1.850 ;
        RECT  0.060 0.660 0.420 0.820 ;
        RECT  1.930 1.100 3.170 1.240 ;
        RECT  1.870 0.710 1.930 1.550 ;
        RECT  1.810 0.710 1.870 1.830 ;
        RECT  1.770 0.710 1.810 0.930 ;
        RECT  1.750 1.430 1.810 1.830 ;
        RECT  3.470 1.420 3.630 1.970 ;
        RECT  3.410 1.420 3.470 1.540 ;
        RECT  3.290 0.710 3.410 1.540 ;
        RECT  3.190 0.710 3.290 0.930 ;
        RECT  4.010 0.420 4.250 0.590 ;
        RECT  3.070 0.470 4.010 0.590 ;
        RECT  2.950 0.470 3.070 0.980 ;
        RECT  2.205 0.860 2.950 0.980 ;
        RECT  2.085 0.470 2.205 0.980 ;
        RECT  1.640 0.470 2.085 0.590 ;
        RECT  1.520 0.470 1.640 0.820 ;
        RECT  1.130 0.700 1.520 0.820 ;
        RECT  0.970 0.700 1.130 1.570 ;
        RECT  0.730 0.700 0.970 0.860 ;
        RECT  5.310 1.170 5.470 2.050 ;
        RECT  4.010 1.930 5.310 2.050 ;
        RECT  3.850 1.120 4.010 2.050 ;
        RECT  3.730 1.120 3.850 1.240 ;
        RECT  6.230 1.080 6.455 1.240 ;
        RECT  6.110 0.680 6.230 1.240 ;
        RECT  5.710 0.680 6.110 0.800 ;
        RECT  5.710 1.780 5.900 1.940 ;
        RECT  5.590 0.680 5.710 1.940 ;
        RECT  5.090 0.680 5.590 0.840 ;
        RECT  5.090 1.650 5.190 1.810 ;
        RECT  4.970 0.680 5.090 1.810 ;
        RECT  3.570 0.760 3.730 1.240 ;
        RECT  4.480 1.220 4.970 1.380 ;
        RECT  3.900 0.810 4.590 0.970 ;
        RECT  0.730 1.410 0.970 1.570 ;
        RECT  2.230 1.380 3.290 1.540 ;
        RECT  1.630 1.670 1.750 1.830 ;
        RECT  2.010 1.670 2.920 1.830 ;
        RECT  0.060 1.690 0.420 1.850 ;
        LAYER M1 ;
        RECT  6.350 0.490 6.455 0.870 ;
        RECT  6.350 1.650 6.455 2.030 ;
    END
END DFCNQD4

MACRO DFCSND1
    CLASS CORE ;
    FOREIGN DFCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.770 1.280 ;
        RECT  3.770 1.005 4.070 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.680 1.440 6.810 1.600 ;
        RECT  6.710 0.420 6.810 0.900 ;
        RECT  6.810 0.420 6.870 1.600 ;
        RECT  6.870 0.780 6.950 1.600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.400 1.960 7.430 2.100 ;
        RECT  7.430 1.390 7.450 2.100 ;
        RECT  7.430 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.590 2.100 ;
        RECT  7.590 1.960 7.620 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.680 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.000 0.300 ;
        RECT  1.000 -0.300 1.220 0.480 ;
        RECT  1.220 -0.300 2.780 0.300 ;
        RECT  2.780 -0.300 3.000 0.560 ;
        RECT  3.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.000 2.820 ;
        RECT  1.000 2.000 1.220 2.820 ;
        RECT  1.220 2.220 2.440 2.820 ;
        RECT  2.440 1.710 2.590 2.820 ;
        RECT  2.590 2.220 3.680 2.820 ;
        RECT  3.680 2.020 3.900 2.820 ;
        RECT  3.900 2.220 4.860 2.820 ;
        RECT  4.860 1.990 5.080 2.820 ;
        RECT  5.080 2.220 5.640 2.820 ;
        RECT  5.640 2.010 5.860 2.820 ;
        RECT  5.860 2.220 6.420 2.820 ;
        RECT  6.420 2.170 6.640 2.820 ;
        RECT  6.640 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.060 0.470 6.180 0.790 ;
        RECT  6.030 1.490 6.430 1.650 ;
        RECT  6.180 0.630 6.430 0.790 ;
        RECT  6.430 0.630 6.550 1.650 ;
        RECT  6.550 1.050 6.690 1.270 ;
        RECT  4.190 0.710 4.310 1.330 ;
        RECT  4.320 1.965 4.350 2.100 ;
        RECT  4.310 1.210 4.350 1.330 ;
        RECT  4.350 1.210 4.470 2.100 ;
        RECT  4.470 1.750 4.540 2.100 ;
        RECT  4.540 1.750 5.010 1.870 ;
        RECT  5.010 1.380 5.130 1.870 ;
        RECT  5.130 1.380 5.510 1.500 ;
        RECT  5.510 1.160 5.670 1.500 ;
        RECT  0.930 1.080 1.130 1.240 ;
        RECT  0.930 0.680 1.530 0.800 ;
        RECT  1.530 0.470 1.650 0.800 ;
        RECT  1.650 0.470 1.910 0.590 ;
        RECT  1.910 0.420 2.110 0.590 ;
        RECT  2.110 0.420 2.130 0.800 ;
        RECT  2.130 0.470 2.230 0.800 ;
        RECT  2.230 0.680 3.120 0.800 ;
        RECT  3.120 0.470 3.240 0.800 ;
        RECT  3.240 0.470 3.930 0.590 ;
        RECT  3.930 0.430 4.150 0.590 ;
        RECT  4.150 0.470 4.540 0.590 ;
        RECT  4.540 0.430 4.760 0.590 ;
        RECT  2.930 1.910 3.340 2.050 ;
        RECT  3.340 1.780 3.460 2.050 ;
        RECT  3.460 1.780 4.040 1.900 ;
        RECT  4.040 1.780 4.200 2.070 ;
        RECT  2.260 0.920 3.370 1.040 ;
        RECT  3.370 0.720 3.490 1.660 ;
        RECT  3.490 0.720 3.920 0.880 ;
        RECT  3.490 1.500 4.160 1.660 ;
        RECT  1.770 0.710 1.800 0.930 ;
        RECT  1.800 0.710 1.920 1.880 ;
        RECT  1.920 0.710 1.940 1.280 ;
        RECT  1.940 1.160 3.030 1.280 ;
        RECT  3.030 1.160 3.250 1.300 ;
        RECT  2.220 1.400 2.800 1.560 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 2.050 ;
        RECT  0.540 1.910 0.620 2.050 ;
        RECT  0.620 1.910 0.860 2.070 ;
        RECT  5.000 0.470 6.060 0.590 ;
        RECT  4.880 0.470 5.000 0.830 ;
        RECT  4.720 0.710 4.880 0.830 ;
        RECT  4.720 1.470 4.850 1.630 ;
        RECT  4.600 0.710 4.720 1.630 ;
        RECT  7.300 1.030 7.330 1.270 ;
        RECT  7.180 1.030 7.300 1.890 ;
        RECT  5.910 1.770 7.180 1.890 ;
        RECT  5.910 1.210 6.140 1.370 ;
        RECT  5.790 0.710 5.910 1.890 ;
        RECT  5.120 0.710 5.790 0.850 ;
        RECT  5.250 1.620 5.790 1.780 ;
        RECT  4.430 0.710 4.600 0.870 ;
        RECT  4.050 0.710 4.190 0.870 ;
        RECT  0.780 0.680 0.930 1.760 ;
        RECT  2.710 1.910 2.930 2.070 ;
        RECT  3.250 1.500 3.370 1.660 ;
        RECT  1.620 1.720 1.800 1.880 ;
        RECT  2.060 1.400 2.220 1.970 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFCSND1

MACRO DFCSND2
    CLASS CORE ;
    FOREIGN DFCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 7.270 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 1.410 7.770 1.810 ;
        RECT  7.660 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.820 1.810 ;
        RECT  7.820 0.780 7.850 1.810 ;
        RECT  7.850 0.780 7.910 1.530 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.320 1.940 8.350 2.100 ;
        RECT  8.350 1.390 8.410 2.100 ;
        RECT  8.350 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.510 2.100 ;
        RECT  8.510 1.940 8.540 2.100 ;
        RECT  8.510 0.780 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.760 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.090 0.300 ;
        RECT  1.090 -0.300 1.310 0.490 ;
        RECT  1.310 -0.300 2.860 0.300 ;
        RECT  2.860 -0.300 3.080 0.560 ;
        RECT  3.080 -0.300 5.050 0.300 ;
        RECT  5.050 -0.300 5.270 0.490 ;
        RECT  5.270 -0.300 7.230 0.300 ;
        RECT  7.230 -0.300 7.450 0.340 ;
        RECT  7.450 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.090 2.820 ;
        RECT  1.090 2.000 1.310 2.820 ;
        RECT  1.310 2.220 2.530 2.820 ;
        RECT  2.530 1.710 2.670 2.820 ;
        RECT  2.670 2.220 3.760 2.820 ;
        RECT  3.760 2.020 3.980 2.820 ;
        RECT  3.980 2.220 4.935 2.820 ;
        RECT  4.935 2.030 5.155 2.820 ;
        RECT  5.155 2.220 6.410 2.820 ;
        RECT  6.410 2.010 6.630 2.820 ;
        RECT  6.630 2.220 7.215 2.820 ;
        RECT  7.215 2.180 7.435 2.820 ;
        RECT  7.435 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.220 0.470 2.310 0.800 ;
        RECT  2.310 0.680 3.200 0.800 ;
        RECT  3.200 0.470 3.320 0.800 ;
        RECT  3.320 0.470 4.010 0.590 ;
        RECT  4.010 0.430 4.230 0.590 ;
        RECT  4.230 0.470 4.620 0.590 ;
        RECT  4.620 0.430 4.860 0.590 ;
        RECT  3.010 1.910 3.420 2.050 ;
        RECT  3.420 1.780 3.540 2.050 ;
        RECT  3.540 1.780 4.150 1.900 ;
        RECT  4.150 1.780 4.310 2.100 ;
        RECT  3.330 1.500 3.450 1.660 ;
        RECT  2.580 0.920 3.450 1.040 ;
        RECT  3.450 0.720 3.570 1.660 ;
        RECT  3.570 0.720 4.000 0.880 ;
        RECT  3.570 1.500 4.240 1.660 ;
        RECT  1.860 0.710 1.880 0.930 ;
        RECT  1.880 0.710 1.920 1.930 ;
        RECT  1.920 0.710 2.000 1.550 ;
        RECT  2.000 0.710 2.020 1.300 ;
        RECT  2.020 1.180 3.110 1.300 ;
        RECT  3.110 1.160 3.330 1.300 ;
        RECT  2.310 1.420 2.880 1.560 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.060 0.720 1.280 ;
        RECT  2.190 0.420 2.220 0.800 ;
        RECT  2.000 0.420 2.190 0.590 ;
        RECT  1.610 0.470 2.000 0.590 ;
        RECT  1.490 0.470 1.610 0.870 ;
        RECT  1.190 0.710 1.490 0.870 ;
        RECT  1.030 0.710 1.190 1.620 ;
        RECT  0.730 0.710 1.030 0.870 ;
        RECT  0.970 1.460 1.030 1.620 ;
        RECT  6.200 1.030 6.360 1.500 ;
        RECT  5.390 1.380 6.200 1.500 ;
        RECT  5.230 1.030 5.390 1.500 ;
        RECT  5.150 1.380 5.230 1.500 ;
        RECT  5.030 1.380 5.150 1.870 ;
        RECT  4.590 1.750 5.030 1.870 ;
        RECT  4.550 1.750 4.590 2.100 ;
        RECT  4.430 1.210 4.550 2.100 ;
        RECT  4.390 1.210 4.430 1.330 ;
        RECT  4.270 0.710 4.390 1.330 ;
        RECT  7.510 1.080 7.650 1.240 ;
        RECT  7.390 0.720 7.510 1.650 ;
        RECT  7.170 0.720 7.390 0.840 ;
        RECT  6.780 1.490 7.390 1.650 ;
        RECT  7.010 0.470 7.170 0.840 ;
        RECT  5.580 0.470 7.010 0.590 ;
        RECT  5.460 0.470 5.580 0.830 ;
        RECT  4.800 0.710 5.460 0.830 ;
        RECT  4.800 1.460 4.910 1.620 ;
        RECT  4.680 0.710 4.800 1.620 ;
        RECT  8.200 1.050 8.290 1.270 ;
        RECT  8.080 1.050 8.200 2.050 ;
        RECT  7.300 1.930 8.080 2.050 ;
        RECT  7.180 1.770 7.300 2.050 ;
        RECT  6.660 1.770 7.180 1.890 ;
        RECT  6.660 1.050 6.690 1.270 ;
        RECT  6.540 0.710 6.660 1.890 ;
        RECT  5.700 0.710 6.540 0.850 ;
        RECT  4.510 0.710 4.680 0.850 ;
        RECT  4.130 0.710 4.270 0.850 ;
        RECT  5.310 1.620 6.540 1.780 ;
        RECT  0.750 1.460 0.970 1.880 ;
        RECT  2.790 1.910 3.010 2.070 ;
        RECT  2.340 0.920 2.580 1.060 ;
        RECT  1.760 1.430 1.880 1.930 ;
        RECT  2.150 1.420 2.310 1.970 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFCSND2

MACRO DFCSND4
    CLASS CORE ;
    FOREIGN DFCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 7.270 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.490 1.600 7.950 1.760 ;
        RECT  7.640 0.490 7.950 0.870 ;
        RECT  7.950 0.490 8.370 1.760 ;
        RECT  8.370 1.600 8.540 1.760 ;
        RECT  8.370 0.490 8.600 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.120 1.650 9.550 2.030 ;
        RECT  9.120 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 2.030 ;
        RECT  9.970 1.650 10.080 2.030 ;
        RECT  9.970 0.490 10.080 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.760 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.095 0.300 ;
        RECT  1.095 -0.300 1.315 0.490 ;
        RECT  1.315 -0.300 2.865 0.300 ;
        RECT  2.865 -0.300 3.085 0.560 ;
        RECT  3.085 -0.300 5.060 0.300 ;
        RECT  5.060 -0.300 5.280 0.590 ;
        RECT  5.280 -0.300 10.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.090 2.820 ;
        RECT  1.090 2.000 1.310 2.820 ;
        RECT  1.310 2.220 2.530 2.820 ;
        RECT  2.530 1.710 2.670 2.820 ;
        RECT  2.670 2.220 2.950 2.820 ;
        RECT  2.950 2.180 3.170 2.820 ;
        RECT  3.170 2.220 3.760 2.820 ;
        RECT  3.760 2.020 3.980 2.820 ;
        RECT  3.980 2.220 4.930 2.820 ;
        RECT  4.930 2.030 5.150 2.820 ;
        RECT  5.150 2.220 6.410 2.820 ;
        RECT  6.410 2.010 6.630 2.820 ;
        RECT  6.630 2.220 8.710 2.820 ;
        RECT  8.710 2.180 8.930 2.820 ;
        RECT  8.930 2.220 10.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.010 1.910 3.420 2.050 ;
        RECT  3.420 1.780 3.540 2.050 ;
        RECT  3.540 1.780 4.150 1.900 ;
        RECT  4.150 1.780 4.310 2.100 ;
        RECT  3.330 1.500 3.450 1.660 ;
        RECT  2.580 0.920 3.450 1.040 ;
        RECT  3.450 0.720 3.570 1.660 ;
        RECT  3.570 0.720 4.000 0.880 ;
        RECT  3.570 1.500 4.240 1.660 ;
        RECT  1.860 0.710 1.880 0.930 ;
        RECT  1.880 0.710 1.920 1.930 ;
        RECT  1.920 0.710 2.000 1.550 ;
        RECT  2.000 0.710 2.020 1.300 ;
        RECT  2.020 1.180 3.110 1.300 ;
        RECT  3.110 1.160 3.330 1.300 ;
        RECT  2.310 1.420 2.880 1.560 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.060 0.720 1.280 ;
        RECT  4.620 0.430 4.860 0.590 ;
        RECT  4.230 0.470 4.620 0.590 ;
        RECT  4.010 0.430 4.230 0.590 ;
        RECT  3.325 0.470 4.010 0.590 ;
        RECT  3.205 0.470 3.325 0.800 ;
        RECT  2.310 0.680 3.205 0.800 ;
        RECT  2.220 0.470 2.310 0.800 ;
        RECT  2.190 0.420 2.220 0.800 ;
        RECT  2.000 0.420 2.190 0.590 ;
        RECT  1.610 0.470 2.000 0.590 ;
        RECT  1.490 0.470 1.610 0.870 ;
        RECT  0.960 0.710 1.490 0.870 ;
        RECT  0.970 1.110 1.205 1.330 ;
        RECT  0.960 1.110 0.970 1.800 ;
        RECT  0.840 0.710 0.960 1.800 ;
        RECT  0.730 0.710 0.840 0.870 ;
        RECT  6.200 1.030 6.360 1.500 ;
        RECT  5.390 1.380 6.200 1.500 ;
        RECT  5.230 1.020 5.390 1.500 ;
        RECT  5.150 1.380 5.230 1.500 ;
        RECT  5.030 1.380 5.150 1.870 ;
        RECT  4.590 1.750 5.030 1.870 ;
        RECT  4.550 1.750 4.590 2.100 ;
        RECT  4.430 1.210 4.550 2.100 ;
        RECT  4.390 1.210 4.430 1.330 ;
        RECT  4.270 0.710 4.390 1.330 ;
        RECT  7.520 1.080 7.640 1.240 ;
        RECT  7.400 0.720 7.520 1.480 ;
        RECT  7.200 0.720 7.400 0.840 ;
        RECT  7.350 1.360 7.400 1.480 ;
        RECT  7.230 1.360 7.350 1.650 ;
        RECT  6.780 1.490 7.230 1.650 ;
        RECT  6.980 0.420 7.200 0.840 ;
        RECT  5.580 0.470 6.980 0.590 ;
        RECT  5.460 0.470 5.580 0.830 ;
        RECT  4.800 0.710 5.460 0.830 ;
        RECT  4.800 1.460 4.910 1.620 ;
        RECT  4.680 0.710 4.800 1.620 ;
        RECT  8.870 1.080 9.240 1.240 ;
        RECT  8.750 1.080 8.870 2.050 ;
        RECT  7.300 1.930 8.750 2.050 ;
        RECT  7.180 1.770 7.300 2.050 ;
        RECT  6.660 1.770 7.180 1.890 ;
        RECT  6.660 1.050 6.690 1.270 ;
        RECT  6.540 0.710 6.660 1.890 ;
        RECT  5.700 0.710 6.540 0.870 ;
        RECT  5.310 1.620 6.540 1.780 ;
        RECT  4.510 0.710 4.680 0.850 ;
        RECT  4.130 0.710 4.270 0.850 ;
        RECT  0.730 1.640 0.840 1.800 ;
        RECT  2.790 1.910 3.010 2.060 ;
        RECT  2.340 0.920 2.580 1.060 ;
        RECT  1.760 1.430 1.880 1.930 ;
        RECT  2.150 1.420 2.310 1.970 ;
        RECT  0.060 1.640 0.420 1.800 ;
        LAYER M1 ;
        RECT  9.120 1.650 9.335 2.030 ;
        RECT  9.120 0.490 9.335 0.870 ;
        RECT  8.585 0.490 8.600 0.870 ;
        RECT  7.640 0.490 7.735 0.870 ;
        RECT  7.490 1.600 7.735 1.760 ;
    END
END DFCSND4

MACRO DFD1
    CLASS CORE ;
    FOREIGN DFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 1.960 5.510 2.100 ;
        RECT  5.510 0.420 5.670 2.100 ;
        RECT  5.670 1.960 5.700 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.960 4.710 2.100 ;
        RECT  4.710 1.390 4.870 2.100 ;
        RECT  4.870 1.390 4.890 1.515 ;
        RECT  4.720 0.710 4.890 0.870 ;
        RECT  4.870 1.960 4.900 2.100 ;
        RECT  4.890 0.710 5.030 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.030 2.820 ;
        RECT  1.030 2.030 1.250 2.820 ;
        RECT  1.250 2.220 2.320 2.820 ;
        RECT  2.320 2.030 2.540 2.820 ;
        RECT  2.540 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.740 1.650 1.210 1.810 ;
        RECT  0.980 0.710 1.210 0.870 ;
        RECT  1.210 0.710 1.370 1.810 ;
        RECT  1.370 0.470 1.510 0.870 ;
        RECT  1.510 0.470 1.910 0.590 ;
        RECT  1.910 0.430 2.130 0.590 ;
        RECT  2.130 0.470 2.970 0.590 ;
        RECT  2.970 0.430 3.190 0.590 ;
        RECT  3.190 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.460 1.290 ;
        RECT  3.460 0.470 3.530 1.560 ;
        RECT  3.530 1.170 3.600 1.560 ;
        RECT  2.700 1.750 2.860 1.910 ;
        RECT  2.410 0.760 2.860 0.920 ;
        RECT  2.860 0.760 2.980 1.910 ;
        RECT  1.710 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  2.070 1.510 2.580 1.630 ;
        RECT  2.580 1.060 2.740 1.630 ;
        RECT  0.070 0.680 0.420 0.840 ;
        RECT  0.420 0.680 0.540 1.795 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  4.230 1.290 4.350 1.450 ;
        RECT  4.110 1.290 4.230 2.050 ;
        RECT  3.290 1.930 4.110 2.050 ;
        RECT  4.600 1.050 4.770 1.270 ;
        RECT  4.590 0.710 4.600 1.270 ;
        RECT  4.510 0.710 4.590 1.730 ;
        RECT  4.470 0.710 4.510 2.090 ;
        RECT  4.100 0.710 4.470 0.850 ;
        RECT  4.350 1.610 4.470 2.090 ;
        RECT  5.240 0.470 5.390 1.290 ;
        RECT  3.810 0.470 5.240 0.590 ;
        RECT  3.810 0.950 3.840 1.810 ;
        RECT  3.720 0.470 3.810 1.810 ;
        RECT  3.650 0.470 3.720 1.050 ;
        RECT  3.560 1.690 3.720 1.810 ;
        RECT  3.960 0.710 4.100 1.160 ;
        RECT  3.130 0.710 3.290 2.050 ;
        RECT  0.760 0.420 0.980 0.870 ;
        RECT  2.250 0.760 2.410 1.320 ;
        RECT  1.720 1.640 1.950 1.800 ;
        RECT  0.070 1.635 0.420 1.795 ;
    END
END DFD1

MACRO DFD2
    CLASS CORE ;
    FOREIGN DFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.060 1.940 6.090 2.100 ;
        RECT  6.090 1.390 6.170 2.100 ;
        RECT  6.090 0.420 6.170 0.900 ;
        RECT  6.170 0.420 6.250 2.100 ;
        RECT  6.250 1.940 6.280 2.100 ;
        RECT  6.250 0.780 6.310 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.350 1.940 5.380 2.100 ;
        RECT  5.380 1.390 5.530 2.100 ;
        RECT  5.330 0.710 5.530 0.870 ;
        RECT  5.530 0.710 5.540 2.100 ;
        RECT  5.540 1.940 5.570 2.100 ;
        RECT  5.540 0.710 5.670 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 4.210 0.300 ;
        RECT  4.210 -0.300 4.430 0.340 ;
        RECT  4.430 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.030 2.820 ;
        RECT  1.030 2.030 1.250 2.820 ;
        RECT  1.250 2.220 2.320 2.820 ;
        RECT  2.320 2.030 2.540 2.820 ;
        RECT  2.540 2.220 4.210 2.820 ;
        RECT  4.210 2.180 4.430 2.820 ;
        RECT  4.430 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.410 0.760 2.835 0.920 ;
        RECT  2.835 0.760 2.960 1.910 ;
        RECT  1.710 0.710 1.990 0.870 ;
        RECT  1.990 0.710 2.110 1.800 ;
        RECT  2.110 1.480 2.120 1.800 ;
        RECT  2.120 1.480 2.570 1.630 ;
        RECT  2.570 1.050 2.715 1.630 ;
        RECT  0.070 0.680 0.420 0.840 ;
        RECT  0.420 0.680 0.540 1.950 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  2.700 1.750 2.835 1.910 ;
        RECT  3.635 1.320 3.690 1.560 ;
        RECT  3.515 0.470 3.635 1.560 ;
        RECT  2.140 0.470 3.515 0.590 ;
        RECT  1.920 0.430 2.140 0.590 ;
        RECT  1.560 0.470 1.920 0.590 ;
        RECT  1.390 0.470 1.560 0.870 ;
        RECT  1.370 0.710 1.390 0.870 ;
        RECT  1.210 0.710 1.370 1.810 ;
        RECT  0.980 0.710 1.210 0.870 ;
        RECT  0.740 1.650 1.210 1.810 ;
        RECT  4.570 1.030 4.730 1.510 ;
        RECT  4.350 1.390 4.570 1.510 ;
        RECT  4.230 1.390 4.350 2.050 ;
        RECT  3.290 1.930 4.230 2.050 ;
        RECT  5.015 1.080 5.410 1.240 ;
        RECT  5.010 0.710 5.015 1.240 ;
        RECT  4.850 0.710 5.010 1.750 ;
        RECT  4.310 0.710 4.850 0.870 ;
        RECT  4.845 1.630 4.850 1.750 ;
        RECT  4.625 1.630 4.845 2.050 ;
        RECT  5.950 1.080 6.050 1.240 ;
        RECT  5.830 0.470 5.950 1.240 ;
        RECT  4.010 0.470 5.830 0.590 ;
        RECT  3.860 0.470 4.010 1.810 ;
        RECT  3.770 1.660 3.860 1.810 ;
        RECT  4.170 0.710 4.310 1.270 ;
        RECT  3.130 0.710 3.290 2.050 ;
        RECT  0.760 0.420 0.980 0.870 ;
        RECT  2.250 0.760 2.410 1.320 ;
        RECT  1.720 1.640 1.990 1.800 ;
        RECT  0.070 1.790 0.420 1.950 ;
    END
END DFD2

MACRO DFD4
    CLASS CORE ;
    FOREIGN DFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.650 7.630 2.030 ;
        RECT  7.290 0.490 7.630 0.870 ;
        RECT  7.630 0.490 8.050 2.030 ;
        RECT  8.050 1.650 8.200 2.030 ;
        RECT  8.050 0.490 8.200 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.910 1.650 6.350 2.030 ;
        RECT  5.890 0.760 6.350 0.920 ;
        RECT  6.350 0.760 6.770 2.030 ;
        RECT  6.770 1.650 6.820 2.030 ;
        RECT  6.770 0.760 6.820 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.300 0.300 ;
        RECT  2.300 -0.300 2.520 0.340 ;
        RECT  2.520 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.030 2.820 ;
        RECT  1.030 2.030 1.250 2.820 ;
        RECT  1.250 2.220 2.320 2.820 ;
        RECT  2.320 2.030 2.540 2.820 ;
        RECT  2.540 2.220 4.820 2.820 ;
        RECT  4.820 2.180 5.040 2.820 ;
        RECT  5.040 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  0.420 0.760 0.540 1.760 ;
        RECT  0.290 0.760 0.420 0.880 ;
        RECT  0.290 1.640 0.420 1.760 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  2.550 1.050 2.710 1.630 ;
        RECT  2.110 1.510 2.550 1.630 ;
        RECT  1.990 0.710 2.110 1.800 ;
        RECT  1.690 0.710 1.990 0.870 ;
        RECT  2.830 0.760 2.950 1.910 ;
        RECT  2.390 0.760 2.830 0.920 ;
        RECT  2.700 1.750 2.830 1.910 ;
        RECT  3.670 1.320 3.700 1.560 ;
        RECT  3.540 0.470 3.670 1.560 ;
        RECT  2.110 0.470 3.540 0.590 ;
        RECT  1.890 0.430 2.110 0.590 ;
        RECT  1.510 0.470 1.890 0.590 ;
        RECT  1.390 0.470 1.510 0.850 ;
        RECT  1.370 0.730 1.390 0.850 ;
        RECT  1.210 0.730 1.370 1.530 ;
        RECT  0.980 0.730 1.210 0.850 ;
        RECT  0.980 1.410 1.210 1.530 ;
        RECT  0.760 0.430 0.980 0.850 ;
        RECT  5.250 1.030 5.410 1.480 ;
        RECT  5.065 1.360 5.250 1.480 ;
        RECT  4.945 1.360 5.065 2.010 ;
        RECT  3.290 1.890 4.945 2.010 ;
        RECT  5.680 1.080 6.020 1.240 ;
        RECT  5.560 0.710 5.680 1.750 ;
        RECT  5.025 0.710 5.560 0.870 ;
        RECT  5.410 1.600 5.560 1.750 ;
        RECT  5.250 1.600 5.410 2.100 ;
        RECT  4.905 0.710 5.025 1.170 ;
        RECT  4.340 1.050 4.905 1.170 ;
        RECT  7.170 1.080 7.400 1.240 ;
        RECT  7.050 0.470 7.170 1.240 ;
        RECT  4.725 0.470 7.050 0.590 ;
        RECT  3.960 1.610 4.745 1.770 ;
        RECT  4.575 0.470 4.725 0.810 ;
        RECT  3.960 0.650 4.575 0.810 ;
        RECT  3.820 0.650 3.960 1.770 ;
        RECT  4.180 1.050 4.340 1.290 ;
        RECT  3.790 0.650 3.820 0.810 ;
        RECT  3.130 0.710 3.290 2.010 ;
        RECT  0.760 1.410 0.980 1.830 ;
        RECT  2.230 0.760 2.390 1.230 ;
        RECT  1.720 1.640 1.990 1.800 ;
        RECT  0.070 1.640 0.290 2.060 ;
        LAYER M1 ;
        RECT  5.890 0.760 6.135 0.920 ;
        RECT  7.290 0.490 7.415 0.870 ;
        RECT  5.910 1.650 6.135 2.030 ;
        RECT  7.290 1.650 7.415 2.030 ;
    END
END DFD4

MACRO DFKCND1
    CLASS CORE ;
    FOREIGN DFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.800 1.940 5.830 2.100 ;
        RECT  5.830 1.390 5.850 2.100 ;
        RECT  5.830 0.420 5.850 0.900 ;
        RECT  5.850 0.420 5.990 2.100 ;
        RECT  5.990 1.940 6.020 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.060 1.860 5.210 2.020 ;
        RECT  5.110 0.710 5.210 0.930 ;
        RECT  5.210 0.710 5.350 2.020 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.650 1.515 ;
        RECT  1.650 1.210 1.810 1.515 ;
        RECT  1.810 1.285 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.710 0.300 ;
        RECT  2.710 -0.300 2.930 0.920 ;
        RECT  2.930 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 4.380 2.820 ;
        RECT  4.380 2.180 4.600 2.820 ;
        RECT  4.600 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.970 1.050 5.090 1.270 ;
        RECT  3.580 0.760 3.700 1.830 ;
        RECT  3.700 1.670 3.770 1.830 ;
        RECT  3.770 1.670 3.890 2.050 ;
        RECT  3.890 1.930 4.570 2.050 ;
        RECT  4.570 1.140 4.690 2.050 ;
        RECT  4.690 1.140 4.730 1.380 ;
        RECT  3.620 0.470 3.820 0.610 ;
        RECT  3.820 0.470 3.940 1.550 ;
        RECT  3.940 1.430 4.080 1.550 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  3.180 0.730 3.340 1.210 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  2.310 0.710 2.430 1.980 ;
        RECT  2.430 1.330 2.470 1.980 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  0.930 1.790 0.950 2.030 ;
        RECT  0.930 0.430 0.950 0.880 ;
        RECT  0.950 0.760 1.420 0.880 ;
        RECT  1.420 0.760 1.540 1.090 ;
        RECT  1.540 0.970 2.030 1.090 ;
        RECT  2.030 0.970 2.190 1.450 ;
        RECT  0.070 0.480 0.510 0.640 ;
        RECT  0.510 0.480 0.670 1.980 ;
        RECT  4.850 0.710 4.970 1.720 ;
        RECT  4.440 0.710 4.850 0.870 ;
        RECT  4.810 1.480 4.850 1.720 ;
        RECT  5.700 1.050 5.730 1.290 ;
        RECT  5.580 0.470 5.700 1.290 ;
        RECT  4.180 0.470 5.580 0.590 ;
        RECT  4.200 1.190 4.320 1.810 ;
        RECT  4.180 1.190 4.200 1.310 ;
        RECT  4.030 1.670 4.200 1.810 ;
        RECT  4.300 0.710 4.440 1.070 ;
        RECT  4.060 0.470 4.180 1.310 ;
        RECT  3.560 0.760 3.580 1.000 ;
        RECT  3.400 0.450 3.620 0.610 ;
        RECT  2.550 1.070 3.180 1.210 ;
        RECT  2.000 0.710 2.310 0.850 ;
        RECT  0.790 0.430 0.930 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.820 0.510 1.980 ;
    END
END DFKCND1

MACRO DFKCND2
    CLASS CORE ;
    FOREIGN DFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.610 1.930 6.640 2.100 ;
        RECT  6.640 1.390 6.800 2.100 ;
        RECT  6.800 1.390 6.810 1.515 ;
        RECT  6.670 0.420 6.810 0.900 ;
        RECT  6.800 1.930 6.830 2.100 ;
        RECT  6.810 0.420 6.840 1.515 ;
        RECT  6.840 0.780 6.950 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.880 1.940 5.910 2.100 ;
        RECT  5.910 1.390 6.070 2.100 ;
        RECT  6.070 1.940 6.100 2.100 ;
        RECT  6.070 1.390 6.130 1.515 ;
        RECT  5.860 0.710 6.130 0.870 ;
        RECT  6.130 0.710 6.310 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.110 1.370 1.315 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.870 ;
        RECT  2.990 -0.300 7.010 0.300 ;
        RECT  7.010 -0.300 7.230 0.340 ;
        RECT  7.230 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 7.010 2.820 ;
        RECT  7.010 2.180 7.230 2.820 ;
        RECT  7.230 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.790 0.430 0.840 0.940 ;
        RECT  0.840 0.430 0.950 2.030 ;
        RECT  0.950 0.760 0.960 2.030 ;
        RECT  0.960 0.760 1.950 0.880 ;
        RECT  1.950 0.760 2.070 1.430 ;
        RECT  2.070 1.210 2.190 1.430 ;
        RECT  0.070 0.690 0.510 0.850 ;
        RECT  0.510 0.690 0.670 1.805 ;
        RECT  0.670 1.090 0.710 1.310 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  2.430 1.330 2.470 1.980 ;
        RECT  2.310 0.680 2.430 1.980 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  3.180 0.710 3.340 1.210 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  4.030 0.450 4.250 0.610 ;
        RECT  3.940 1.430 4.100 1.550 ;
        RECT  3.940 0.470 4.030 0.610 ;
        RECT  5.060 1.050 5.300 1.270 ;
        RECT  4.940 1.050 5.060 2.050 ;
        RECT  3.890 1.930 4.940 2.050 ;
        RECT  3.770 1.670 3.890 2.050 ;
        RECT  3.700 1.670 3.770 1.830 ;
        RECT  3.580 0.490 3.700 1.830 ;
        RECT  5.600 1.050 5.990 1.270 ;
        RECT  5.480 0.710 5.600 1.620 ;
        RECT  4.770 0.710 5.480 0.870 ;
        RECT  5.340 1.500 5.480 1.620 ;
        RECT  5.180 1.500 5.340 2.000 ;
        RECT  6.550 1.080 6.680 1.240 ;
        RECT  6.430 0.470 6.550 1.240 ;
        RECT  4.500 0.470 6.430 0.590 ;
        RECT  4.500 1.670 4.660 1.810 ;
        RECT  4.380 0.470 4.500 1.810 ;
        RECT  4.230 0.830 4.380 0.950 ;
        RECT  4.030 1.670 4.380 1.810 ;
        RECT  4.620 0.710 4.770 1.290 ;
        RECT  4.060 0.730 4.230 0.950 ;
        RECT  3.560 0.490 3.580 1.000 ;
        RECT  3.820 0.470 3.940 1.550 ;
        RECT  2.630 1.070 3.180 1.210 ;
        RECT  2.190 0.680 2.310 0.900 ;
        RECT  0.790 1.500 0.840 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.645 0.510 1.805 ;
    END
END DFKCND2

MACRO DFKCND4
    CLASS CORE ;
    FOREIGN DFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 1.650 7.950 2.030 ;
        RECT  7.630 0.490 7.950 0.870 ;
        RECT  7.950 0.490 8.370 2.030 ;
        RECT  8.370 1.650 8.540 2.030 ;
        RECT  8.370 0.490 8.540 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.200 1.650 6.670 2.030 ;
        RECT  6.180 0.760 6.670 0.920 ;
        RECT  6.670 0.760 7.090 2.030 ;
        RECT  7.090 1.650 7.150 2.030 ;
        RECT  7.090 0.760 7.170 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.210 1.690 1.430 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.110 1.370 1.315 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.870 ;
        RECT  2.990 -0.300 4.320 0.300 ;
        RECT  4.320 -0.300 4.540 0.340 ;
        RECT  4.540 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 4.340 2.820 ;
        RECT  4.340 2.180 4.560 2.820 ;
        RECT  4.560 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.720 0.510 0.880 ;
        RECT  0.510 0.720 0.670 1.810 ;
        RECT  0.670 1.090 0.710 1.310 ;
        RECT  0.290 1.650 0.510 1.810 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  2.070 1.210 2.190 1.430 ;
        RECT  1.950 0.760 2.070 1.430 ;
        RECT  0.960 0.760 1.950 0.880 ;
        RECT  0.950 0.760 0.960 2.030 ;
        RECT  0.840 0.430 0.950 2.030 ;
        RECT  0.790 0.430 0.840 0.940 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  2.430 1.330 2.470 1.930 ;
        RECT  2.310 0.680 2.430 1.930 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  3.180 0.710 3.340 1.210 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  4.030 0.450 4.250 0.610 ;
        RECT  3.940 1.410 4.100 1.550 ;
        RECT  3.940 0.470 4.030 0.610 ;
        RECT  5.380 1.050 5.620 1.270 ;
        RECT  5.260 1.050 5.380 2.050 ;
        RECT  3.890 1.930 5.260 2.050 ;
        RECT  3.770 1.670 3.890 2.050 ;
        RECT  3.700 1.670 3.770 1.830 ;
        RECT  3.580 0.490 3.700 1.830 ;
        RECT  5.920 1.050 6.240 1.270 ;
        RECT  5.800 0.710 5.920 1.680 ;
        RECT  4.940 0.710 5.800 0.870 ;
        RECT  5.660 1.560 5.800 1.680 ;
        RECT  5.500 1.560 5.660 2.060 ;
        RECT  7.490 1.080 7.735 1.240 ;
        RECT  7.370 0.470 7.490 1.240 ;
        RECT  4.940 0.470 7.370 0.590 ;
        RECT  4.595 1.670 4.980 1.810 ;
        RECT  4.760 0.450 4.940 0.590 ;
        RECT  4.595 0.470 4.760 0.590 ;
        RECT  4.475 0.470 4.595 1.810 ;
        RECT  4.230 0.830 4.475 0.950 ;
        RECT  4.030 1.670 4.475 1.810 ;
        RECT  4.780 0.710 4.940 1.290 ;
        RECT  4.060 0.730 4.230 0.950 ;
        RECT  3.560 0.490 3.580 1.000 ;
        RECT  3.820 0.470 3.940 1.550 ;
        RECT  2.630 1.070 3.180 1.210 ;
        RECT  2.190 0.680 2.310 0.900 ;
        RECT  0.790 1.500 0.840 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.650 0.290 2.070 ;
        LAYER M1 ;
        RECT  7.630 1.650 7.735 2.030 ;
        RECT  7.630 0.490 7.735 0.870 ;
        RECT  6.200 1.650 6.455 2.030 ;
        RECT  6.180 0.760 6.455 0.920 ;
    END
END DFKCND4

MACRO DFKCNQD1
    CLASS CORE ;
    FOREIGN DFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.940 5.150 2.100 ;
        RECT  5.150 1.390 5.210 2.100 ;
        RECT  5.150 0.420 5.210 0.900 ;
        RECT  5.210 0.420 5.310 2.100 ;
        RECT  5.310 1.940 5.340 2.100 ;
        RECT  5.310 0.780 5.350 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.650 1.515 ;
        RECT  1.650 1.210 1.810 1.515 ;
        RECT  1.810 1.285 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.710 0.300 ;
        RECT  2.710 -0.300 2.930 0.920 ;
        RECT  2.930 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 4.380 2.820 ;
        RECT  4.380 2.180 4.600 2.820 ;
        RECT  4.600 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.310 0.710 2.430 1.980 ;
        RECT  2.430 1.330 2.470 1.980 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  0.930 1.790 0.950 2.030 ;
        RECT  0.930 0.430 0.950 0.880 ;
        RECT  0.950 0.760 1.420 0.880 ;
        RECT  1.420 0.760 1.540 1.090 ;
        RECT  1.540 0.970 2.030 1.090 ;
        RECT  2.030 0.970 2.190 1.450 ;
        RECT  0.070 0.480 0.510 0.640 ;
        RECT  0.510 0.480 0.670 1.980 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  3.180 0.730 3.340 1.210 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  3.940 1.430 4.080 1.550 ;
        RECT  3.820 0.470 3.940 1.550 ;
        RECT  3.620 0.470 3.820 0.610 ;
        RECT  4.200 1.190 4.320 1.810 ;
        RECT  4.180 1.190 4.200 1.310 ;
        RECT  4.030 1.670 4.200 1.810 ;
        RECT  4.690 1.140 4.730 1.380 ;
        RECT  4.570 1.140 4.690 2.050 ;
        RECT  3.890 1.930 4.570 2.050 ;
        RECT  3.770 1.670 3.890 2.050 ;
        RECT  3.700 1.670 3.770 1.830 ;
        RECT  3.580 0.760 3.700 1.830 ;
        RECT  4.990 1.050 5.090 1.270 ;
        RECT  4.970 0.570 4.990 1.270 ;
        RECT  4.850 0.570 4.970 1.780 ;
        RECT  4.440 0.570 4.850 0.730 ;
        RECT  4.810 1.540 4.850 1.780 ;
        RECT  3.560 0.760 3.580 1.000 ;
        RECT  4.060 0.560 4.180 1.310 ;
        RECT  3.400 0.450 3.620 0.610 ;
        RECT  2.550 1.070 3.180 1.210 ;
        RECT  2.000 0.710 2.310 0.850 ;
        RECT  0.790 0.430 0.930 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.820 0.510 1.980 ;
        RECT  4.300 0.570 4.440 1.070 ;
    END
END DFKCNQD1

MACRO DFKCNQD2
    CLASS CORE ;
    FOREIGN DFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.630 1.950 5.660 2.090 ;
        RECT  5.660 1.380 5.820 2.090 ;
        RECT  5.820 1.950 5.850 2.090 ;
        RECT  5.820 1.380 5.850 1.515 ;
        RECT  5.630 0.500 5.850 0.920 ;
        RECT  5.850 0.760 5.990 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.110 1.370 1.315 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.870 ;
        RECT  2.990 -0.300 4.410 0.300 ;
        RECT  4.410 -0.300 4.630 0.340 ;
        RECT  4.630 -0.300 5.220 0.300 ;
        RECT  5.220 -0.300 5.440 0.340 ;
        RECT  5.440 -0.300 6.040 0.300 ;
        RECT  6.040 -0.300 6.260 0.340 ;
        RECT  6.260 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 4.410 2.820 ;
        RECT  4.410 2.180 4.630 2.820 ;
        RECT  4.630 2.220 5.220 2.820 ;
        RECT  5.220 2.180 5.440 2.820 ;
        RECT  5.440 2.220 6.040 2.820 ;
        RECT  6.040 2.180 6.260 2.820 ;
        RECT  6.260 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.670 1.090 0.710 1.310 ;
        RECT  0.510 0.690 0.670 1.805 ;
        RECT  0.070 0.690 0.510 0.850 ;
        RECT  2.070 1.210 2.190 1.430 ;
        RECT  1.950 0.760 2.070 1.430 ;
        RECT  0.960 0.760 1.950 0.880 ;
        RECT  0.950 0.760 0.960 2.030 ;
        RECT  0.840 0.430 0.950 2.030 ;
        RECT  0.790 0.430 0.840 0.940 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  2.430 1.330 2.470 1.930 ;
        RECT  2.310 0.680 2.430 1.930 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  3.180 0.710 3.340 1.210 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  3.940 1.410 4.080 1.570 ;
        RECT  3.820 0.450 3.940 1.570 ;
        RECT  4.720 1.080 5.010 1.240 ;
        RECT  4.600 1.080 4.720 1.850 ;
        RECT  3.700 1.690 4.600 1.850 ;
        RECT  3.580 0.750 3.700 1.850 ;
        RECT  5.260 1.080 5.720 1.240 ;
        RECT  5.140 0.710 5.260 1.550 ;
        RECT  4.430 0.710 5.140 0.870 ;
        RECT  5.000 1.430 5.140 1.550 ;
        RECT  4.840 1.430 5.000 1.930 ;
        RECT  4.310 0.710 4.430 1.570 ;
        RECT  3.560 0.750 3.580 1.000 ;
        RECT  3.690 0.450 3.820 0.610 ;
        RECT  2.630 1.070 3.180 1.210 ;
        RECT  2.190 0.680 2.310 0.900 ;
        RECT  0.790 1.500 0.840 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.645 0.510 1.805 ;
        RECT  4.210 1.410 4.310 1.570 ;
    END
END DFKCNQD2

MACRO DFKCNQD4
    CLASS CORE ;
    FOREIGN DFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.540 1.650 6.030 2.030 ;
        RECT  5.540 0.490 6.030 0.870 ;
        RECT  6.030 0.490 6.450 2.030 ;
        RECT  6.450 1.650 6.490 2.030 ;
        RECT  6.450 0.490 6.490 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.110 1.370 1.315 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.120 0.300 ;
        RECT  1.120 -0.300 1.340 0.640 ;
        RECT  1.340 -0.300 2.770 0.300 ;
        RECT  2.770 -0.300 2.990 0.870 ;
        RECT  2.990 -0.300 4.410 0.300 ;
        RECT  4.410 -0.300 4.630 0.340 ;
        RECT  4.630 -0.300 6.680 0.300 ;
        RECT  6.680 -0.300 6.900 0.340 ;
        RECT  6.900 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 1.950 1.730 2.820 ;
        RECT  1.730 2.220 2.910 2.820 ;
        RECT  2.910 1.770 3.130 2.820 ;
        RECT  3.130 2.220 4.410 2.820 ;
        RECT  4.410 2.180 4.630 2.820 ;
        RECT  4.630 2.220 6.680 2.820 ;
        RECT  6.680 2.180 6.900 2.820 ;
        RECT  6.900 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.950 0.760 0.960 2.030 ;
        RECT  0.960 0.760 1.950 0.880 ;
        RECT  1.950 0.760 2.070 1.430 ;
        RECT  2.070 1.210 2.190 1.430 ;
        RECT  0.070 0.480 0.510 0.640 ;
        RECT  0.840 0.430 0.950 2.030 ;
        RECT  0.790 0.430 0.840 0.940 ;
        RECT  2.470 1.330 3.220 1.470 ;
        RECT  2.430 1.330 2.470 1.980 ;
        RECT  2.310 0.680 2.430 1.980 ;
        RECT  2.190 0.680 2.310 0.900 ;
        RECT  0.510 0.480 0.670 1.980 ;
        RECT  0.670 1.090 0.710 1.310 ;
        RECT  3.340 1.090 3.460 1.880 ;
        RECT  3.180 0.710 3.340 1.210 ;
        RECT  3.320 1.640 3.340 1.880 ;
        RECT  3.940 1.410 4.080 1.570 ;
        RECT  3.820 0.450 3.940 1.570 ;
        RECT  4.720 1.080 5.010 1.240 ;
        RECT  4.600 1.080 4.720 1.850 ;
        RECT  3.700 1.690 4.600 1.850 ;
        RECT  3.580 0.750 3.700 1.850 ;
        RECT  5.260 1.080 5.815 1.240 ;
        RECT  5.140 0.750 5.260 1.500 ;
        RECT  5.030 0.750 5.140 0.910 ;
        RECT  5.000 1.380 5.140 1.500 ;
        RECT  4.810 0.490 5.030 0.910 ;
        RECT  5.000 1.950 5.030 2.090 ;
        RECT  4.840 1.380 5.000 2.090 ;
        RECT  4.810 1.950 4.840 2.090 ;
        RECT  4.430 0.750 4.810 0.910 ;
        RECT  4.310 0.750 4.430 1.570 ;
        RECT  4.210 1.410 4.310 1.570 ;
        RECT  3.560 0.750 3.580 1.000 ;
        RECT  3.690 0.450 3.820 0.610 ;
        RECT  2.630 1.070 3.180 1.210 ;
        RECT  0.790 1.500 0.840 2.030 ;
        RECT  1.100 1.670 2.140 1.830 ;
        RECT  0.070 1.820 0.510 1.980 ;
        LAYER M1 ;
        RECT  5.540 1.650 5.815 2.030 ;
        RECT  5.540 0.490 5.815 0.870 ;
    END
END DFKCNQD4

MACRO DFKCSND1
    CLASS CORE ;
    FOREIGN DFKCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.940 6.790 2.100 ;
        RECT  6.790 1.390 6.810 2.100 ;
        RECT  6.790 0.420 6.810 0.900 ;
        RECT  6.810 0.420 6.950 2.100 ;
        RECT  6.950 1.940 6.980 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.940 6.070 2.100 ;
        RECT  6.070 1.390 6.170 2.100 ;
        RECT  6.020 0.710 6.170 0.870 ;
        RECT  6.170 0.710 6.230 2.100 ;
        RECT  6.230 1.940 6.260 2.100 ;
        RECT  6.230 0.710 6.310 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.440 1.650 ;
        RECT  0.870 0.930 1.440 1.050 ;
        RECT  1.440 0.930 1.560 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.110 0.300 ;
        RECT  2.110 -0.300 2.330 0.340 ;
        RECT  2.330 -0.300 3.710 0.300 ;
        RECT  3.710 -0.300 3.930 0.480 ;
        RECT  3.930 -0.300 5.370 0.300 ;
        RECT  5.370 -0.300 5.590 0.340 ;
        RECT  5.590 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.420 2.820 ;
        RECT  1.420 2.180 1.640 2.820 ;
        RECT  1.640 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 3.660 2.820 ;
        RECT  3.660 2.040 3.880 2.820 ;
        RECT  3.880 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.660 1.050 6.690 1.290 ;
        RECT  5.400 1.090 5.710 1.210 ;
        RECT  5.710 0.710 5.870 1.980 ;
        RECT  5.870 1.080 6.050 1.240 ;
        RECT  4.530 0.720 4.660 0.940 ;
        RECT  4.530 1.870 5.410 2.030 ;
        RECT  5.410 1.330 5.530 2.030 ;
        RECT  5.530 1.330 5.570 1.570 ;
        RECT  4.650 1.120 4.780 1.750 ;
        RECT  4.580 0.470 4.780 0.590 ;
        RECT  4.780 0.470 4.810 1.750 ;
        RECT  4.810 0.470 4.900 1.240 ;
        RECT  4.040 1.680 4.170 1.840 ;
        RECT  4.140 0.700 4.170 1.170 ;
        RECT  4.170 0.700 4.290 1.840 ;
        RECT  3.100 0.630 3.230 0.790 ;
        RECT  3.230 0.630 3.350 1.770 ;
        RECT  3.350 1.400 3.890 1.520 ;
        RECT  3.890 1.300 4.050 1.520 ;
        RECT  2.380 0.710 2.510 0.870 ;
        RECT  2.510 0.710 2.630 1.690 ;
        RECT  2.630 1.300 3.070 1.460 ;
        RECT  1.260 0.470 2.770 0.590 ;
        RECT  2.770 0.470 2.930 0.750 ;
        RECT  1.240 1.930 2.770 2.050 ;
        RECT  2.770 1.630 2.930 2.050 ;
        RECT  1.690 0.710 2.020 0.870 ;
        RECT  2.020 0.710 2.140 1.780 ;
        RECT  2.140 1.040 2.380 1.270 ;
        RECT  0.070 0.590 0.350 0.750 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.320 1.310 ;
        RECT  6.540 0.470 6.660 1.290 ;
        RECT  5.160 0.470 6.540 0.590 ;
        RECT  5.140 0.470 5.160 0.890 ;
        RECT  5.020 0.470 5.140 1.750 ;
        RECT  5.260 0.970 5.400 1.210 ;
        RECT  4.930 1.530 5.020 1.750 ;
        RECT  4.410 0.720 4.530 2.030 ;
        RECT  4.360 0.430 4.580 0.590 ;
        RECT  3.600 1.010 4.140 1.170 ;
        RECT  3.100 1.610 3.230 1.770 ;
        RECT  2.380 1.530 2.510 1.690 ;
        RECT  1.100 0.470 1.260 0.810 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  1.690 1.640 2.020 1.780 ;
        RECT  0.070 1.850 0.350 2.010 ;
    END
END DFKCSND1

MACRO DFKCSND2
    CLASS CORE ;
    FOREIGN DFKCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.345 1.950 7.375 2.090 ;
        RECT  7.375 1.380 7.535 2.090 ;
        RECT  7.535 1.950 7.565 2.090 ;
        RECT  7.345 0.500 7.565 0.920 ;
        RECT  7.535 1.380 7.770 1.515 ;
        RECT  7.565 0.800 7.770 0.920 ;
        RECT  7.770 0.800 7.910 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.655 1.960 6.685 2.100 ;
        RECT  6.685 1.390 6.810 2.100 ;
        RECT  6.635 0.760 6.810 0.920 ;
        RECT  6.810 0.760 6.845 2.100 ;
        RECT  6.845 1.960 6.875 2.100 ;
        RECT  6.845 0.760 6.950 1.525 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.440 1.650 ;
        RECT  0.870 0.930 1.440 1.050 ;
        RECT  1.440 0.930 1.560 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.000 0.300 ;
        RECT  2.000 -0.300 2.220 0.340 ;
        RECT  2.220 -0.300 3.670 0.300 ;
        RECT  3.670 -0.300 3.890 0.480 ;
        RECT  3.890 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.420 2.820 ;
        RECT  1.420 2.180 1.640 2.820 ;
        RECT  1.640 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 3.660 2.820 ;
        RECT  3.660 2.040 3.880 2.820 ;
        RECT  3.880 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.170 0.680 4.250 1.840 ;
        RECT  4.250 1.010 4.290 1.840 ;
        RECT  3.100 0.600 3.230 0.760 ;
        RECT  3.230 0.600 3.350 1.770 ;
        RECT  3.350 1.300 4.050 1.520 ;
        RECT  2.380 0.750 2.510 0.910 ;
        RECT  2.510 0.750 2.630 1.690 ;
        RECT  2.630 1.300 3.110 1.460 ;
        RECT  1.260 0.470 2.980 0.620 ;
        RECT  1.240 1.930 2.770 2.050 ;
        RECT  2.770 1.630 2.930 2.050 ;
        RECT  1.690 0.740 2.020 0.885 ;
        RECT  2.020 0.740 2.140 1.795 ;
        RECT  2.140 1.040 2.380 1.270 ;
        RECT  0.070 0.590 0.350 0.750 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.320 1.310 ;
        RECT  4.100 0.680 4.170 1.170 ;
        RECT  4.040 1.680 4.170 1.840 ;
        RECT  4.860 0.430 5.140 0.590 ;
        RECT  4.810 0.430 4.860 1.240 ;
        RECT  4.740 0.430 4.810 1.750 ;
        RECT  5.880 1.080 6.145 1.245 ;
        RECT  5.760 1.080 5.880 2.030 ;
        RECT  4.530 1.870 5.760 2.030 ;
        RECT  4.530 0.730 4.620 0.950 ;
        RECT  6.385 1.050 6.690 1.270 ;
        RECT  6.265 0.750 6.385 1.500 ;
        RECT  5.640 0.750 6.265 0.910 ;
        RECT  6.155 1.380 6.265 1.500 ;
        RECT  6.000 1.380 6.155 1.880 ;
        RECT  5.500 0.750 5.640 1.230 ;
        RECT  7.225 1.080 7.520 1.240 ;
        RECT  7.105 0.470 7.225 1.240 ;
        RECT  5.380 0.470 7.105 0.630 ;
        RECT  5.120 1.590 5.515 1.750 ;
        RECT  5.260 0.470 5.380 0.890 ;
        RECT  5.120 0.720 5.260 0.890 ;
        RECT  4.980 0.720 5.120 1.750 ;
        RECT  5.480 0.990 5.500 1.230 ;
        RECT  4.410 0.730 4.530 2.030 ;
        RECT  4.650 1.120 4.740 1.750 ;
        RECT  3.580 1.010 4.100 1.170 ;
        RECT  3.100 1.610 3.230 1.770 ;
        RECT  2.380 1.530 2.510 1.690 ;
        RECT  1.100 0.470 1.260 0.810 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  1.690 1.635 2.020 1.795 ;
        RECT  0.070 1.850 0.350 2.010 ;
        RECT  4.930 1.530 4.980 1.750 ;
    END
END DFKCSND2

MACRO DFKCSND4
    CLASS CORE ;
    FOREIGN DFKCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.490 1.630 8.910 2.010 ;
        RECT  8.490 0.510 8.910 0.890 ;
        RECT  8.910 0.510 9.330 2.010 ;
        RECT  9.330 1.630 9.460 2.010 ;
        RECT  9.330 0.510 9.460 0.890 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.030 1.630 7.310 2.010 ;
        RECT  7.010 0.760 7.310 0.920 ;
        RECT  7.310 0.760 7.730 2.010 ;
        RECT  7.730 1.630 7.980 2.010 ;
        RECT  7.730 0.760 8.000 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.440 1.650 ;
        RECT  0.870 0.930 1.440 1.050 ;
        RECT  1.440 0.930 1.560 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.670 0.300 ;
        RECT  3.670 -0.300 3.890 0.480 ;
        RECT  3.890 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.420 2.820 ;
        RECT  1.420 2.180 1.640 2.820 ;
        RECT  1.640 2.220 3.660 2.820 ;
        RECT  3.660 2.040 3.880 2.820 ;
        RECT  3.880 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.320 1.310 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.070 0.590 0.350 0.750 ;
        RECT  2.140 1.040 2.380 1.270 ;
        RECT  2.020 0.710 2.140 1.795 ;
        RECT  1.690 0.710 2.020 0.870 ;
        RECT  2.770 1.630 2.930 2.050 ;
        RECT  1.240 1.930 2.770 2.050 ;
        RECT  2.770 0.470 2.930 0.750 ;
        RECT  1.260 0.470 2.770 0.590 ;
        RECT  2.630 1.300 3.070 1.460 ;
        RECT  2.510 0.710 2.630 1.690 ;
        RECT  2.380 0.710 2.510 0.870 ;
        RECT  3.910 1.300 4.050 1.520 ;
        RECT  3.350 1.400 3.910 1.520 ;
        RECT  3.230 0.600 3.350 1.770 ;
        RECT  3.120 0.600 3.230 0.790 ;
        RECT  4.250 1.010 4.290 1.840 ;
        RECT  4.170 0.680 4.250 1.840 ;
        RECT  4.100 0.680 4.170 1.170 ;
        RECT  4.040 1.680 4.170 1.840 ;
        RECT  4.860 0.430 5.140 0.590 ;
        RECT  4.810 0.430 4.860 1.240 ;
        RECT  4.740 0.430 4.810 1.750 ;
        RECT  6.090 1.080 6.410 1.240 ;
        RECT  5.970 1.080 6.090 2.030 ;
        RECT  4.530 1.870 5.970 2.030 ;
        RECT  4.530 0.750 4.620 0.970 ;
        RECT  6.735 1.050 7.090 1.270 ;
        RECT  6.615 0.750 6.735 1.500 ;
        RECT  5.740 0.750 6.615 0.910 ;
        RECT  6.490 1.380 6.615 1.500 ;
        RECT  6.490 1.950 6.520 2.090 ;
        RECT  6.330 1.380 6.490 2.090 ;
        RECT  6.300 1.950 6.330 2.090 ;
        RECT  8.310 1.080 8.600 1.240 ;
        RECT  8.190 0.470 8.310 1.240 ;
        RECT  5.400 0.470 8.190 0.630 ;
        RECT  5.100 1.610 5.810 1.750 ;
        RECT  5.260 0.470 5.400 0.930 ;
        RECT  5.100 0.740 5.260 0.930 ;
        RECT  4.980 0.740 5.100 1.750 ;
        RECT  5.580 0.750 5.740 1.230 ;
        RECT  4.930 1.530 4.980 1.750 ;
        RECT  4.410 0.750 4.530 2.030 ;
        RECT  4.650 1.120 4.740 1.750 ;
        RECT  3.580 1.010 4.100 1.170 ;
        RECT  3.100 1.610 3.230 1.770 ;
        RECT  2.380 1.530 2.510 1.690 ;
        RECT  1.100 0.470 1.260 0.810 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  1.690 1.635 2.020 1.795 ;
        RECT  0.070 1.850 0.350 2.010 ;
        LAYER M1 ;
        RECT  7.945 0.760 8.000 0.920 ;
        RECT  7.010 0.760 7.095 0.920 ;
        RECT  8.490 1.630 8.695 2.010 ;
        RECT  7.945 1.630 7.980 2.010 ;
        RECT  7.030 1.630 7.095 2.010 ;
        RECT  8.490 0.510 8.695 0.890 ;
    END
END DFKCSND4

MACRO DFKSND1
    CLASS CORE ;
    FOREIGN DFKSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.285 1.510 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 1.940 6.470 2.100 ;
        RECT  6.470 1.390 6.490 2.100 ;
        RECT  6.470 0.420 6.490 0.900 ;
        RECT  6.490 0.420 6.630 2.100 ;
        RECT  6.630 1.940 6.660 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.730 1.940 5.760 2.100 ;
        RECT  5.760 1.390 5.850 2.100 ;
        RECT  5.710 0.710 5.850 0.870 ;
        RECT  5.850 0.710 5.920 2.100 ;
        RECT  5.920 1.940 5.950 2.100 ;
        RECT  5.920 0.710 5.990 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.990 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.310 0.300 ;
        RECT  1.310 -0.300 1.530 0.340 ;
        RECT  1.530 -0.300 2.110 0.300 ;
        RECT  2.110 -0.300 2.330 0.340 ;
        RECT  2.330 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.850 ;
        RECT  3.630 -0.300 4.990 0.300 ;
        RECT  4.990 -0.300 5.210 0.340 ;
        RECT  5.210 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 3.480 2.820 ;
        RECT  3.480 1.830 3.700 2.820 ;
        RECT  3.700 2.220 4.990 2.820 ;
        RECT  4.990 2.180 5.210 2.820 ;
        RECT  5.210 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.470 4.850 1.670 ;
        RECT  4.850 0.470 4.870 0.900 ;
        RECT  4.850 1.450 4.890 1.670 ;
        RECT  4.870 0.470 6.230 0.590 ;
        RECT  6.230 0.470 6.350 1.290 ;
        RECT  6.350 1.050 6.370 1.290 ;
        RECT  5.110 1.150 5.420 1.270 ;
        RECT  5.420 0.710 5.580 1.670 ;
        RECT  5.580 1.050 5.730 1.270 ;
        RECT  4.370 1.790 5.290 1.950 ;
        RECT  5.290 1.790 5.450 2.080 ;
        RECT  4.290 0.470 4.490 0.590 ;
        RECT  4.490 0.470 4.610 1.670 ;
        RECT  3.500 1.550 3.990 1.710 ;
        RECT  3.800 0.710 3.990 0.850 ;
        RECT  3.990 0.710 4.110 1.710 ;
        RECT  2.750 0.780 3.040 0.940 ;
        RECT  3.040 0.780 3.160 1.770 ;
        RECT  3.160 0.970 3.680 1.090 ;
        RECT  3.680 0.970 3.840 1.380 ;
        RECT  0.060 0.470 0.420 0.630 ;
        RECT  0.420 0.470 0.540 2.050 ;
        RECT  0.540 1.010 0.660 1.230 ;
        RECT  0.540 1.930 2.510 2.050 ;
        RECT  2.510 1.030 2.670 2.050 ;
        RECT  2.670 1.930 2.960 2.050 ;
        RECT  2.960 1.930 3.200 2.090 ;
        RECT  0.900 1.590 0.940 1.810 ;
        RECT  0.900 0.420 0.940 0.640 ;
        RECT  0.940 0.470 2.910 0.590 ;
        RECT  2.910 0.430 3.150 0.590 ;
        RECT  1.690 0.710 2.270 0.870 ;
        RECT  2.270 0.710 2.390 1.800 ;
        RECT  2.390 0.710 2.590 0.870 ;
        RECT  1.090 1.650 1.640 1.810 ;
        RECT  1.200 1.040 1.640 1.160 ;
        RECT  1.640 1.040 1.800 1.810 ;
        RECT  4.970 1.030 5.110 1.270 ;
        RECT  4.230 0.710 4.370 1.950 ;
        RECT  4.050 0.430 4.290 0.590 ;
        RECT  3.340 1.210 3.500 1.710 ;
        RECT  2.810 1.610 3.040 1.770 ;
        RECT  0.060 1.650 0.420 1.810 ;
        RECT  0.780 0.420 0.900 1.810 ;
        RECT  2.140 1.640 2.270 1.800 ;
        RECT  1.040 0.760 1.200 1.160 ;
    END
END DFKSND1

MACRO DFKSND2
    CLASS CORE ;
    FOREIGN DFKSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.285 1.510 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 1.940 7.070 2.100 ;
        RECT  7.070 1.390 7.130 2.100 ;
        RECT  7.070 0.420 7.130 0.900 ;
        RECT  7.130 0.420 7.230 2.100 ;
        RECT  7.230 1.940 7.260 2.100 ;
        RECT  7.230 0.780 7.270 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.940 6.380 2.100 ;
        RECT  6.380 1.390 6.490 2.100 ;
        RECT  6.330 0.710 6.490 0.870 ;
        RECT  6.490 0.710 6.540 2.100 ;
        RECT  6.540 1.940 6.570 2.100 ;
        RECT  6.540 0.710 6.630 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.990 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.310 0.300 ;
        RECT  1.310 -0.300 1.530 0.340 ;
        RECT  1.530 -0.300 2.000 0.300 ;
        RECT  2.000 -0.300 2.220 0.340 ;
        RECT  2.220 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.850 ;
        RECT  3.630 -0.300 5.080 0.300 ;
        RECT  5.080 -0.300 5.300 0.340 ;
        RECT  5.300 -0.300 5.950 0.300 ;
        RECT  5.950 -0.300 6.170 0.340 ;
        RECT  6.170 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 3.480 2.820 ;
        RECT  3.480 1.830 3.700 2.820 ;
        RECT  3.700 2.220 5.100 2.820 ;
        RECT  5.100 2.180 5.320 2.820 ;
        RECT  5.320 2.220 5.950 2.820 ;
        RECT  5.950 2.180 6.170 2.820 ;
        RECT  6.170 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.780 3.040 0.940 ;
        RECT  3.040 0.780 3.160 1.770 ;
        RECT  3.160 0.970 3.680 1.090 ;
        RECT  3.680 0.970 3.840 1.380 ;
        RECT  0.060 0.470 0.420 0.630 ;
        RECT  0.420 0.470 0.540 2.050 ;
        RECT  0.540 1.010 0.660 1.230 ;
        RECT  0.540 1.930 2.510 2.050 ;
        RECT  2.510 1.030 2.650 2.050 ;
        RECT  2.650 1.030 2.670 1.220 ;
        RECT  2.650 1.930 2.960 2.050 ;
        RECT  2.960 1.930 3.200 2.100 ;
        RECT  0.900 1.590 0.940 1.810 ;
        RECT  0.900 0.420 0.940 0.640 ;
        RECT  0.940 0.470 2.910 0.590 ;
        RECT  2.910 0.430 3.150 0.590 ;
        RECT  1.690 0.710 2.270 0.870 ;
        RECT  2.270 0.710 2.390 1.810 ;
        RECT  2.390 0.710 2.590 0.870 ;
        RECT  1.090 1.650 1.640 1.810 ;
        RECT  1.200 1.040 1.640 1.160 ;
        RECT  1.640 1.040 1.800 1.810 ;
        RECT  3.990 0.710 4.110 1.710 ;
        RECT  3.800 0.710 3.990 0.850 ;
        RECT  3.500 1.550 3.990 1.710 ;
        RECT  4.490 0.470 4.610 1.700 ;
        RECT  4.290 0.470 4.490 0.590 ;
        RECT  5.440 1.050 5.540 1.270 ;
        RECT  5.320 1.050 5.440 1.510 ;
        RECT  5.130 1.390 5.320 1.510 ;
        RECT  5.010 1.390 5.130 2.050 ;
        RECT  4.370 1.890 5.010 2.050 ;
        RECT  5.820 1.080 6.370 1.240 ;
        RECT  5.700 0.710 5.820 1.780 ;
        RECT  5.090 0.710 5.700 0.870 ;
        RECT  5.500 1.620 5.700 1.780 ;
        RECT  6.950 1.050 7.010 1.270 ;
        RECT  6.830 0.470 6.950 1.270 ;
        RECT  4.850 0.470 6.830 0.590 ;
        RECT  4.850 1.550 4.890 1.770 ;
        RECT  4.730 0.470 4.850 1.770 ;
        RECT  4.970 0.710 5.090 1.270 ;
        RECT  4.230 0.720 4.370 2.050 ;
        RECT  4.050 0.420 4.290 0.590 ;
        RECT  3.340 1.210 3.500 1.710 ;
        RECT  2.770 1.610 3.040 1.770 ;
        RECT  0.060 1.650 0.420 1.810 ;
        RECT  0.780 0.420 0.900 1.810 ;
        RECT  2.140 1.650 2.270 1.810 ;
        RECT  1.040 0.760 1.200 1.160 ;
    END
END DFKSND2

MACRO DFKSND4
    CLASS CORE ;
    FOREIGN DFKSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.280 1.370 1.515 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.650 8.590 2.030 ;
        RECT  8.270 0.490 8.590 0.870 ;
        RECT  8.590 0.490 9.010 2.030 ;
        RECT  9.010 1.650 9.180 2.030 ;
        RECT  9.010 0.490 9.180 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.890 1.650 7.310 2.030 ;
        RECT  6.870 0.750 7.310 0.910 ;
        RECT  7.310 0.750 7.730 2.030 ;
        RECT  7.730 1.650 7.800 2.030 ;
        RECT  7.730 0.750 7.820 0.910 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.990 2.470 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 1.480 0.300 ;
        RECT  1.480 -0.300 1.700 0.340 ;
        RECT  1.700 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.340 ;
        RECT  2.390 -0.300 3.580 0.300 ;
        RECT  3.580 -0.300 3.800 0.850 ;
        RECT  3.800 -0.300 5.090 0.300 ;
        RECT  5.090 -0.300 5.310 0.340 ;
        RECT  5.310 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.180 0.670 2.820 ;
        RECT  0.670 2.220 1.680 2.820 ;
        RECT  1.680 2.180 1.900 2.820 ;
        RECT  1.900 2.220 3.650 2.820 ;
        RECT  3.650 1.830 3.870 2.820 ;
        RECT  3.870 2.220 5.110 2.820 ;
        RECT  5.110 2.180 5.330 2.820 ;
        RECT  5.330 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.820 1.030 2.840 1.220 ;
        RECT  2.820 1.930 3.130 2.050 ;
        RECT  3.130 1.930 3.370 2.100 ;
        RECT  1.060 0.470 3.080 0.590 ;
        RECT  3.080 0.430 3.320 0.590 ;
        RECT  2.060 0.710 2.180 1.810 ;
        RECT  2.180 1.650 2.560 1.810 ;
        RECT  2.180 0.710 2.760 0.870 ;
        RECT  1.640 0.725 1.760 1.160 ;
        RECT  1.260 1.650 1.780 1.810 ;
        RECT  1.760 1.040 1.780 1.160 ;
        RECT  1.780 1.040 1.940 1.810 ;
        RECT  2.680 1.030 2.820 2.050 ;
        RECT  0.630 1.930 2.680 2.050 ;
        RECT  0.630 1.050 0.720 1.270 ;
        RECT  0.510 0.725 0.630 2.050 ;
        RECT  0.280 0.725 0.510 0.885 ;
        RECT  0.280 1.930 0.510 2.050 ;
        RECT  0.060 0.465 0.280 0.885 ;
        RECT  3.850 0.970 4.010 1.380 ;
        RECT  3.330 0.970 3.850 1.090 ;
        RECT  3.210 0.780 3.330 1.770 ;
        RECT  2.920 0.780 3.210 0.940 ;
        RECT  4.150 0.690 4.270 1.710 ;
        RECT  3.950 0.690 4.150 0.850 ;
        RECT  3.670 1.550 4.150 1.710 ;
        RECT  6.015 1.080 6.270 1.240 ;
        RECT  5.895 1.080 6.015 2.050 ;
        RECT  4.540 1.890 5.895 2.050 ;
        RECT  6.520 1.080 7.055 1.240 ;
        RECT  6.400 0.750 6.520 1.500 ;
        RECT  6.390 1.950 6.420 2.090 ;
        RECT  5.675 0.750 6.400 0.910 ;
        RECT  6.390 1.380 6.400 1.500 ;
        RECT  6.230 1.380 6.390 2.090 ;
        RECT  6.200 1.950 6.230 2.090 ;
        RECT  8.150 1.080 8.375 1.240 ;
        RECT  8.030 0.470 8.150 1.240 ;
        RECT  4.970 0.470 8.030 0.630 ;
        RECT  4.970 1.530 5.750 1.690 ;
        RECT  4.850 0.470 4.970 1.690 ;
        RECT  4.710 0.760 4.850 0.920 ;
        RECT  5.515 0.750 5.675 1.290 ;
        RECT  4.390 0.700 4.540 2.050 ;
        RECT  3.510 1.210 3.670 1.710 ;
        RECT  2.940 1.610 3.210 1.770 ;
        RECT  0.060 1.635 0.280 2.050 ;
        RECT  0.840 0.470 1.060 1.810 ;
        RECT  1.880 0.710 2.060 0.870 ;
        RECT  1.180 0.725 1.640 0.885 ;
        LAYER M1 ;
        RECT  8.270 1.650 8.375 2.030 ;
        RECT  8.270 0.490 8.375 0.870 ;
        RECT  6.890 1.650 7.095 2.030 ;
        RECT  6.870 0.750 7.095 0.910 ;
    END
END DFKSND4

MACRO DFNCND1
    CLASS CORE ;
    FOREIGN DFNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.940 6.790 2.100 ;
        RECT  6.790 0.420 6.950 2.100 ;
        RECT  6.950 1.940 6.980 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.920 1.940 5.950 2.100 ;
        RECT  5.950 1.390 6.110 2.100 ;
        RECT  6.110 1.940 6.140 2.100 ;
        RECT  6.110 1.390 6.170 1.515 ;
        RECT  5.900 0.710 6.170 0.830 ;
        RECT  6.170 0.710 6.310 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.660 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.285 4.910 1.515 ;
        RECT  4.910 1.190 5.070 1.515 ;
        RECT  5.070 1.285 5.350 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.000 0.300 ;
        RECT  1.000 -0.300 1.220 0.480 ;
        RECT  1.220 -0.300 2.660 0.300 ;
        RECT  2.660 -0.300 2.820 0.740 ;
        RECT  2.820 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.940 0.550 ;
        RECT  4.940 -0.300 6.340 0.300 ;
        RECT  6.340 -0.300 6.560 0.340 ;
        RECT  6.560 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.000 2.820 ;
        RECT  1.000 2.000 1.220 2.820 ;
        RECT  1.220 2.220 2.420 2.820 ;
        RECT  2.420 2.030 2.640 2.820 ;
        RECT  2.640 2.220 3.050 2.820 ;
        RECT  3.050 1.670 3.270 2.820 ;
        RECT  3.270 2.220 4.610 2.820 ;
        RECT  4.610 2.180 4.830 2.820 ;
        RECT  4.830 2.220 5.440 2.820 ;
        RECT  5.440 2.180 5.660 2.820 ;
        RECT  5.660 2.220 6.340 2.820 ;
        RECT  6.340 2.180 6.560 2.820 ;
        RECT  6.560 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.730 0.950 5.390 1.070 ;
        RECT  5.390 0.710 5.550 1.070 ;
        RECT  5.550 0.950 5.890 1.070 ;
        RECT  5.890 0.950 6.050 1.270 ;
        RECT  3.720 1.120 3.840 1.240 ;
        RECT  3.840 1.120 4.000 2.050 ;
        RECT  4.000 1.930 5.470 2.050 ;
        RECT  5.470 1.190 5.630 2.050 ;
        RECT  2.070 0.430 2.190 0.980 ;
        RECT  2.190 0.860 2.940 0.980 ;
        RECT  2.940 0.470 3.060 0.980 ;
        RECT  3.060 0.470 4.020 0.590 ;
        RECT  4.020 0.430 4.240 0.590 ;
        RECT  3.180 0.710 3.280 0.930 ;
        RECT  3.280 0.710 3.400 1.540 ;
        RECT  3.400 1.420 3.460 1.540 ;
        RECT  3.460 1.420 3.620 1.990 ;
        RECT  1.780 0.710 1.900 1.800 ;
        RECT  1.900 0.710 1.930 1.260 ;
        RECT  1.930 1.100 3.160 1.260 ;
        RECT  2.240 1.670 2.670 1.800 ;
        RECT  2.670 1.670 2.910 1.830 ;
        RECT  0.940 1.050 1.050 1.270 ;
        RECT  0.940 1.645 1.400 1.765 ;
        RECT  1.400 1.645 1.520 2.050 ;
        RECT  1.520 1.920 2.060 2.050 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 2.050 ;
        RECT  0.540 1.910 0.620 2.050 ;
        RECT  0.620 1.910 0.860 2.070 ;
        RECT  4.730 1.650 5.270 1.810 ;
        RECT  6.510 0.470 6.670 1.290 ;
        RECT  5.240 0.470 6.510 0.590 ;
        RECT  5.120 0.470 5.240 0.830 ;
        RECT  4.450 0.670 5.120 0.830 ;
        RECT  4.330 0.670 4.450 1.810 ;
        RECT  3.890 0.830 4.330 0.990 ;
        RECT  4.570 0.950 4.730 1.810 ;
        RECT  3.560 0.770 3.720 1.240 ;
        RECT  1.900 0.430 2.070 0.590 ;
        RECT  2.220 1.380 3.280 1.540 ;
        RECT  1.640 1.640 1.780 1.800 ;
        RECT  2.020 1.660 2.240 1.800 ;
        RECT  0.780 0.660 0.940 1.765 ;
        RECT  0.060 1.640 0.420 1.800 ;
        RECT  4.180 1.650 4.330 1.810 ;
    END
END DFNCND1

MACRO DFNCND2
    CLASS CORE ;
    FOREIGN DFNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.350 1.940 7.380 2.100 ;
        RECT  7.380 1.390 7.450 2.100 ;
        RECT  7.380 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.540 2.100 ;
        RECT  7.540 1.940 7.570 2.100 ;
        RECT  7.540 0.780 7.590 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.560 1.940 6.590 2.100 ;
        RECT  6.590 1.390 6.750 2.100 ;
        RECT  6.750 1.940 6.780 2.100 ;
        RECT  6.750 1.390 6.810 1.515 ;
        RECT  6.560 0.710 6.810 0.830 ;
        RECT  6.810 0.710 6.950 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.750 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.960 1.125 6.120 1.625 ;
        RECT  6.120 1.465 6.170 1.625 ;
        RECT  6.170 1.465 6.310 2.075 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.020 0.300 ;
        RECT  1.020 -0.300 1.240 0.490 ;
        RECT  1.240 -0.300 2.730 0.300 ;
        RECT  2.730 -0.300 2.890 0.570 ;
        RECT  2.890 -0.300 4.790 0.300 ;
        RECT  4.790 -0.300 5.010 0.550 ;
        RECT  5.010 -0.300 6.120 0.300 ;
        RECT  6.120 -0.300 6.340 0.340 ;
        RECT  6.340 -0.300 6.955 0.300 ;
        RECT  6.955 -0.300 7.175 0.340 ;
        RECT  7.175 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.010 2.820 ;
        RECT  1.010 2.000 1.230 2.820 ;
        RECT  1.230 2.220 2.490 2.820 ;
        RECT  2.490 2.030 2.710 2.820 ;
        RECT  2.710 2.220 3.120 2.820 ;
        RECT  3.120 1.670 3.340 2.820 ;
        RECT  3.340 2.220 4.675 2.820 ;
        RECT  4.675 2.180 4.910 2.820 ;
        RECT  4.910 2.220 6.955 2.820 ;
        RECT  6.955 2.180 7.175 2.820 ;
        RECT  7.175 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 0.690 3.010 0.810 ;
        RECT  3.010 0.470 3.130 0.810 ;
        RECT  3.130 0.470 4.090 0.590 ;
        RECT  4.090 0.430 4.310 0.590 ;
        RECT  3.250 0.710 3.350 0.930 ;
        RECT  3.350 0.710 3.470 1.470 ;
        RECT  3.470 1.350 3.530 1.470 ;
        RECT  3.530 1.350 3.690 1.990 ;
        RECT  1.780 1.390 1.870 1.800 ;
        RECT  1.840 0.710 1.870 0.930 ;
        RECT  1.870 0.710 1.900 1.800 ;
        RECT  1.900 0.710 1.990 1.510 ;
        RECT  1.990 0.710 2.000 1.190 ;
        RECT  2.000 1.050 3.230 1.190 ;
        RECT  0.780 0.680 0.840 0.900 ;
        RECT  0.840 0.680 0.980 1.760 ;
        RECT  0.980 0.950 0.990 1.760 ;
        RECT  0.990 0.950 1.250 1.110 ;
        RECT  0.990 1.640 1.370 1.760 ;
        RECT  1.370 1.640 1.490 2.050 ;
        RECT  1.490 1.930 2.200 2.050 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.050 0.720 1.270 ;
        RECT  2.140 0.430 2.260 0.810 ;
        RECT  5.440 1.190 5.560 2.050 ;
        RECT  5.340 1.190 5.440 1.390 ;
        RECT  4.070 1.930 5.440 2.050 ;
        RECT  3.910 1.090 4.070 2.050 ;
        RECT  3.800 1.090 3.910 1.210 ;
        RECT  6.440 0.950 6.600 1.270 ;
        RECT  6.320 0.755 6.440 1.070 ;
        RECT  5.800 0.755 6.320 0.875 ;
        RECT  5.800 1.775 6.030 1.935 ;
        RECT  5.680 0.755 5.800 1.935 ;
        RECT  5.620 0.755 5.680 1.070 ;
        RECT  5.460 0.710 5.620 1.070 ;
        RECT  4.800 0.950 5.460 1.070 ;
        RECT  4.800 1.650 5.320 1.810 ;
        RECT  7.260 1.050 7.300 1.290 ;
        RECT  7.140 0.470 7.260 1.290 ;
        RECT  5.310 0.470 7.140 0.590 ;
        RECT  5.190 0.470 5.310 0.830 ;
        RECT  4.520 0.670 5.190 0.830 ;
        RECT  4.400 0.670 4.520 1.810 ;
        RECT  3.970 0.810 4.400 0.970 ;
        RECT  4.250 1.650 4.400 1.810 ;
        RECT  4.640 0.950 4.800 1.810 ;
        RECT  3.640 0.760 3.800 1.210 ;
        RECT  1.970 0.430 2.140 0.590 ;
        RECT  2.290 1.310 3.350 1.470 ;
        RECT  1.740 1.560 1.780 1.800 ;
        RECT  2.070 1.600 2.980 1.760 ;
        RECT  0.780 1.540 0.840 1.760 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFNCND2

MACRO DFNCND4
    CLASS CORE ;
    FOREIGN DFNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.590 1.650 8.910 2.030 ;
        RECT  8.590 0.490 8.910 0.870 ;
        RECT  8.910 0.490 9.330 2.030 ;
        RECT  9.330 1.650 9.500 2.030 ;
        RECT  9.330 0.490 9.500 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.210 1.650 7.310 2.030 ;
        RECT  7.210 0.760 7.310 0.920 ;
        RECT  7.310 0.760 7.730 2.030 ;
        RECT  7.730 1.650 8.120 2.030 ;
        RECT  7.730 0.760 8.140 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.005 1.700 1.225 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.980 1.190 6.140 1.445 ;
        RECT  6.140 1.285 6.170 1.445 ;
        RECT  6.170 1.285 6.310 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.020 0.300 ;
        RECT  1.020 -0.300 1.240 0.480 ;
        RECT  1.240 -0.300 2.730 0.300 ;
        RECT  2.730 -0.300 2.890 0.620 ;
        RECT  2.890 -0.300 4.790 0.300 ;
        RECT  4.790 -0.300 5.010 0.550 ;
        RECT  5.010 -0.300 6.080 0.300 ;
        RECT  6.080 -0.300 6.300 0.340 ;
        RECT  6.300 -0.300 6.820 0.300 ;
        RECT  6.820 -0.300 7.040 0.340 ;
        RECT  7.040 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.020 2.820 ;
        RECT  1.020 2.000 1.240 2.820 ;
        RECT  1.240 2.220 3.060 2.820 ;
        RECT  3.060 2.025 3.290 2.820 ;
        RECT  3.290 2.220 4.670 2.820 ;
        RECT  4.670 2.180 4.910 2.820 ;
        RECT  4.910 2.220 6.210 2.820 ;
        RECT  6.210 2.180 6.430 2.820 ;
        RECT  6.430 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.050 0.720 1.270 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  1.480 1.930 2.185 2.050 ;
        RECT  1.360 1.635 1.480 2.050 ;
        RECT  1.240 1.635 1.360 1.755 ;
        RECT  1.080 0.710 1.240 1.755 ;
        RECT  0.730 0.710 1.080 0.870 ;
        RECT  2.000 1.040 3.200 1.170 ;
        RECT  1.970 0.710 2.000 1.170 ;
        RECT  1.840 0.710 1.970 1.730 ;
        RECT  3.540 1.330 3.700 1.990 ;
        RECT  3.470 1.330 3.540 1.450 ;
        RECT  3.350 0.710 3.470 1.450 ;
        RECT  3.250 0.710 3.350 0.930 ;
        RECT  2.440 1.330 3.350 1.450 ;
        RECT  4.090 0.430 4.310 0.590 ;
        RECT  3.130 0.470 4.090 0.590 ;
        RECT  3.010 0.470 3.130 0.860 ;
        RECT  2.260 0.740 3.010 0.860 ;
        RECT  2.140 0.430 2.260 0.860 ;
        RECT  5.440 1.190 5.560 2.050 ;
        RECT  5.400 1.190 5.440 1.410 ;
        RECT  4.080 1.930 5.440 2.050 ;
        RECT  3.920 1.090 4.080 2.050 ;
        RECT  3.800 1.090 3.920 1.210 ;
        RECT  6.690 0.950 6.850 1.290 ;
        RECT  5.800 0.950 6.690 1.070 ;
        RECT  5.800 1.760 6.050 1.920 ;
        RECT  5.680 0.950 5.800 1.920 ;
        RECT  5.620 0.950 5.680 1.070 ;
        RECT  5.460 0.750 5.620 1.070 ;
        RECT  4.800 0.950 5.460 1.070 ;
        RECT  4.800 1.650 5.320 1.810 ;
        RECT  8.470 1.080 8.695 1.240 ;
        RECT  8.350 0.470 8.470 1.240 ;
        RECT  7.090 0.470 8.350 0.590 ;
        RECT  6.970 0.470 7.090 1.650 ;
        RECT  5.310 0.470 6.970 0.630 ;
        RECT  6.500 1.490 6.970 1.650 ;
        RECT  5.190 0.470 5.310 0.830 ;
        RECT  4.520 0.670 5.190 0.830 ;
        RECT  4.400 0.670 4.520 1.690 ;
        RECT  3.970 0.810 4.400 0.970 ;
        RECT  4.640 0.950 4.800 1.810 ;
        RECT  3.640 0.760 3.800 1.210 ;
        RECT  4.250 1.530 4.400 1.690 ;
        RECT  1.970 0.430 2.140 0.590 ;
        RECT  2.200 1.290 2.440 1.450 ;
        RECT  1.700 1.570 1.840 1.730 ;
        RECT  2.100 1.610 3.030 1.770 ;
        RECT  0.730 1.595 1.080 1.755 ;
        RECT  0.060 1.640 0.420 1.800 ;
        LAYER M1 ;
        RECT  7.945 0.760 8.140 0.920 ;
        RECT  7.945 1.650 8.120 2.030 ;
        RECT  8.590 0.490 8.695 0.870 ;
        RECT  8.590 1.650 8.695 2.030 ;
    END
END DFNCND4

MACRO DFNCSND1
    CLASS CORE ;
    FOREIGN DFNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.770 1.280 ;
        RECT  3.770 1.005 4.070 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.680 1.440 6.810 1.600 ;
        RECT  6.710 0.420 6.810 0.900 ;
        RECT  6.810 0.420 6.870 1.600 ;
        RECT  6.870 0.780 6.950 1.600 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.400 1.960 7.430 2.100 ;
        RECT  7.430 1.390 7.450 2.100 ;
        RECT  7.430 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.590 2.100 ;
        RECT  7.590 1.960 7.620 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.660 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.000 0.300 ;
        RECT  1.000 -0.300 1.220 0.480 ;
        RECT  1.220 -0.300 2.780 0.300 ;
        RECT  2.780 -0.300 3.000 0.560 ;
        RECT  3.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.000 2.820 ;
        RECT  1.000 2.000 1.220 2.820 ;
        RECT  1.220 2.220 2.460 2.820 ;
        RECT  2.460 1.710 2.600 2.820 ;
        RECT  2.600 2.220 3.680 2.820 ;
        RECT  3.680 2.020 3.900 2.820 ;
        RECT  3.900 2.220 4.860 2.820 ;
        RECT  4.860 1.990 5.080 2.820 ;
        RECT  5.080 2.220 5.640 2.820 ;
        RECT  5.640 2.010 5.860 2.820 ;
        RECT  5.860 2.220 6.420 2.820 ;
        RECT  6.420 2.170 6.640 2.820 ;
        RECT  6.640 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.880 0.470 5.000 0.830 ;
        RECT  5.000 0.470 6.060 0.590 ;
        RECT  6.060 0.470 6.180 0.790 ;
        RECT  6.030 1.490 6.430 1.650 ;
        RECT  6.180 0.630 6.430 0.790 ;
        RECT  6.430 0.630 6.550 1.650 ;
        RECT  6.550 1.050 6.690 1.270 ;
        RECT  4.190 0.710 4.310 1.330 ;
        RECT  4.320 1.960 4.350 2.100 ;
        RECT  4.310 1.210 4.350 1.330 ;
        RECT  4.350 1.210 4.470 2.100 ;
        RECT  4.470 1.750 4.540 2.100 ;
        RECT  4.540 1.750 5.010 1.870 ;
        RECT  5.010 1.380 5.130 1.870 ;
        RECT  5.130 1.380 5.510 1.500 ;
        RECT  5.510 1.160 5.670 1.500 ;
        RECT  2.180 0.680 3.120 0.800 ;
        RECT  3.120 0.470 3.240 0.800 ;
        RECT  3.240 0.470 3.930 0.590 ;
        RECT  3.930 0.430 4.150 0.590 ;
        RECT  4.150 0.470 4.540 0.590 ;
        RECT  4.540 0.430 4.760 0.590 ;
        RECT  2.900 1.880 3.340 2.020 ;
        RECT  3.340 1.780 3.460 2.020 ;
        RECT  3.460 1.780 4.040 1.900 ;
        RECT  4.040 1.780 4.200 2.070 ;
        RECT  3.250 1.500 3.370 1.660 ;
        RECT  2.530 0.920 3.370 1.040 ;
        RECT  3.370 0.720 3.490 1.660 ;
        RECT  3.490 0.720 3.920 0.880 ;
        RECT  3.490 1.500 4.160 1.660 ;
        RECT  1.780 0.450 1.900 1.780 ;
        RECT  1.900 0.450 1.920 1.300 ;
        RECT  1.920 1.180 3.030 1.300 ;
        RECT  3.030 1.160 3.250 1.300 ;
        RECT  2.150 1.420 2.270 1.840 ;
        RECT  2.270 1.420 2.800 1.560 ;
        RECT  0.940 1.080 1.130 1.240 ;
        RECT  0.940 1.635 1.375 1.755 ;
        RECT  1.375 1.635 1.495 2.050 ;
        RECT  1.495 1.930 1.800 2.050 ;
        RECT  1.800 1.930 1.950 2.100 ;
        RECT  1.950 1.960 2.060 2.100 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 2.050 ;
        RECT  0.540 1.910 0.620 2.050 ;
        RECT  0.620 1.910 0.860 2.070 ;
        RECT  4.720 0.710 4.880 0.830 ;
        RECT  4.720 1.470 4.850 1.630 ;
        RECT  4.600 0.710 4.720 1.630 ;
        RECT  7.300 1.030 7.330 1.270 ;
        RECT  7.180 1.030 7.300 1.890 ;
        RECT  5.910 1.770 7.180 1.890 ;
        RECT  5.910 1.210 6.140 1.370 ;
        RECT  5.790 0.710 5.910 1.890 ;
        RECT  5.120 0.710 5.790 0.850 ;
        RECT  4.430 0.710 4.600 0.870 ;
        RECT  4.050 0.710 4.190 0.870 ;
        RECT  2.040 0.680 2.180 1.040 ;
        RECT  2.740 1.880 2.900 2.100 ;
        RECT  2.310 0.920 2.530 1.060 ;
        RECT  1.620 1.620 1.780 1.780 ;
        RECT  5.250 1.620 5.790 1.780 ;
        RECT  2.030 1.680 2.150 1.840 ;
        RECT  0.780 0.660 0.940 1.755 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFNCSND1

MACRO DFNCSND2
    CLASS CORE ;
    FOREIGN DFNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.070 1.015 7.130 1.235 ;
        RECT  7.130 0.725 7.270 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.630 1.410 7.770 1.810 ;
        RECT  7.660 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.820 1.810 ;
        RECT  7.820 0.780 7.850 1.810 ;
        RECT  7.850 0.780 7.910 1.530 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.320 1.940 8.350 2.100 ;
        RECT  8.350 1.390 8.410 2.100 ;
        RECT  8.350 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.510 2.100 ;
        RECT  8.510 1.940 8.540 2.100 ;
        RECT  8.510 0.780 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.030 1.770 1.250 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.090 0.300 ;
        RECT  1.090 -0.300 1.310 0.490 ;
        RECT  1.310 -0.300 3.070 0.300 ;
        RECT  3.070 -0.300 3.290 0.530 ;
        RECT  3.290 -0.300 5.140 0.300 ;
        RECT  5.140 -0.300 5.360 0.490 ;
        RECT  5.360 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.090 2.820 ;
        RECT  1.090 2.000 1.320 2.820 ;
        RECT  1.320 2.220 2.620 2.820 ;
        RECT  2.620 1.710 2.760 2.820 ;
        RECT  2.760 2.220 3.850 2.820 ;
        RECT  3.850 2.020 4.070 2.820 ;
        RECT  4.070 2.220 5.020 2.820 ;
        RECT  5.020 2.030 5.240 2.820 ;
        RECT  5.240 2.220 6.500 2.820 ;
        RECT  6.500 2.010 6.720 2.820 ;
        RECT  6.720 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.100 1.910 3.510 2.050 ;
        RECT  3.510 1.780 3.630 2.050 ;
        RECT  3.630 1.780 4.210 1.900 ;
        RECT  4.210 1.780 4.370 2.100 ;
        RECT  2.550 0.890 3.650 1.010 ;
        RECT  3.650 0.720 3.770 1.660 ;
        RECT  3.770 0.720 4.090 0.880 ;
        RECT  3.770 1.500 4.330 1.660 ;
        RECT  1.930 0.450 2.070 1.745 ;
        RECT  2.070 0.450 2.090 1.250 ;
        RECT  2.090 1.130 3.310 1.250 ;
        RECT  3.310 1.130 3.530 1.310 ;
        RECT  2.390 1.400 2.990 1.560 ;
        RECT  0.730 0.710 0.840 0.870 ;
        RECT  0.840 0.710 0.970 1.800 ;
        RECT  0.970 1.050 1.065 1.270 ;
        RECT  0.970 1.680 1.500 1.800 ;
        RECT  1.500 1.680 1.630 2.050 ;
        RECT  1.630 1.930 1.980 2.050 ;
        RECT  1.980 1.930 2.200 2.070 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.060 0.720 1.280 ;
        RECT  4.710 0.430 4.950 0.590 ;
        RECT  4.320 0.470 4.710 0.590 ;
        RECT  4.100 0.430 4.320 0.590 ;
        RECT  3.530 0.470 4.100 0.590 ;
        RECT  3.410 0.470 3.530 0.770 ;
        RECT  2.370 0.650 3.410 0.770 ;
        RECT  6.290 1.030 6.450 1.500 ;
        RECT  5.410 1.380 6.290 1.500 ;
        RECT  5.250 1.030 5.410 1.500 ;
        RECT  5.240 1.380 5.250 1.500 ;
        RECT  5.120 1.380 5.240 1.870 ;
        RECT  4.710 1.750 5.120 1.870 ;
        RECT  4.610 1.750 4.710 2.100 ;
        RECT  4.490 1.210 4.610 2.100 ;
        RECT  4.480 1.210 4.490 1.330 ;
        RECT  4.360 0.710 4.480 1.330 ;
        RECT  7.510 1.080 7.650 1.240 ;
        RECT  7.390 0.470 7.510 1.650 ;
        RECT  7.210 0.470 7.390 0.590 ;
        RECT  6.870 1.490 7.390 1.650 ;
        RECT  6.990 0.430 7.210 0.590 ;
        RECT  5.640 0.470 6.990 0.590 ;
        RECT  5.520 0.470 5.640 0.830 ;
        RECT  4.890 0.710 5.520 0.830 ;
        RECT  4.890 1.460 5.000 1.620 ;
        RECT  4.770 0.710 4.890 1.620 ;
        RECT  8.200 1.050 8.290 1.270 ;
        RECT  8.080 1.050 8.200 2.050 ;
        RECT  7.140 1.930 8.080 2.050 ;
        RECT  7.020 1.770 7.140 2.050 ;
        RECT  6.730 1.770 7.020 1.890 ;
        RECT  6.730 1.155 6.760 1.375 ;
        RECT  6.720 1.155 6.730 1.890 ;
        RECT  6.610 0.710 6.720 1.890 ;
        RECT  6.600 0.710 6.610 1.780 ;
        RECT  5.770 0.710 6.600 0.850 ;
        RECT  4.600 0.710 4.770 0.850 ;
        RECT  4.220 0.710 4.360 0.850 ;
        RECT  2.210 0.650 2.370 0.960 ;
        RECT  2.880 1.910 3.100 2.070 ;
        RECT  3.420 1.500 3.650 1.660 ;
        RECT  1.780 1.585 1.930 1.745 ;
        RECT  2.230 1.400 2.390 1.810 ;
        RECT  0.730 1.640 0.840 1.800 ;
        RECT  0.060 1.640 0.420 1.800 ;
        RECT  5.400 1.620 6.600 1.780 ;
    END
END DFNCSND2

MACRO DFNCSND4
    CLASS CORE ;
    FOREIGN DFNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.010 1.075 7.130 1.235 ;
        RECT  7.130 0.725 7.270 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.570 1.600 7.950 1.760 ;
        RECT  7.720 0.490 7.950 0.870 ;
        RECT  7.950 0.490 8.370 1.760 ;
        RECT  8.370 1.600 8.580 1.760 ;
        RECT  8.370 0.490 8.640 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.160 1.650 9.550 2.030 ;
        RECT  9.160 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 2.030 ;
        RECT  9.970 1.650 10.080 2.030 ;
        RECT  9.970 0.490 10.080 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.775 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.090 0.300 ;
        RECT  1.090 -0.300 1.310 0.490 ;
        RECT  1.310 -0.300 3.060 0.300 ;
        RECT  3.060 -0.300 3.280 0.490 ;
        RECT  3.280 -0.300 5.130 0.300 ;
        RECT  5.130 -0.300 5.350 0.490 ;
        RECT  5.350 -0.300 10.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.090 2.820 ;
        RECT  1.090 2.000 1.310 2.820 ;
        RECT  1.310 2.220 2.640 2.820 ;
        RECT  2.640 1.700 2.760 2.820 ;
        RECT  2.760 2.220 3.840 2.820 ;
        RECT  3.840 2.020 4.060 2.820 ;
        RECT  4.060 2.220 5.010 2.820 ;
        RECT  5.010 2.030 5.230 2.820 ;
        RECT  5.230 2.220 6.490 2.820 ;
        RECT  6.490 2.010 6.710 2.820 ;
        RECT  6.710 2.220 8.750 2.820 ;
        RECT  8.750 2.180 8.970 2.820 ;
        RECT  8.970 2.220 10.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.700 0.430 4.940 0.590 ;
        RECT  3.110 1.910 3.500 2.050 ;
        RECT  3.500 1.780 3.620 2.050 ;
        RECT  3.620 1.780 4.230 1.900 ;
        RECT  4.230 1.780 4.390 2.100 ;
        RECT  2.540 0.850 3.640 0.970 ;
        RECT  3.640 0.720 3.760 1.660 ;
        RECT  3.760 0.720 4.080 0.880 ;
        RECT  3.760 1.500 4.320 1.660 ;
        RECT  1.940 0.450 2.060 1.650 ;
        RECT  2.060 0.450 2.100 1.270 ;
        RECT  2.100 1.150 3.300 1.270 ;
        RECT  3.300 1.150 3.520 1.290 ;
        RECT  2.290 1.400 2.410 1.810 ;
        RECT  2.410 1.400 2.960 1.560 ;
        RECT  0.750 0.450 0.850 0.870 ;
        RECT  0.850 0.450 0.970 2.060 ;
        RECT  0.970 1.050 1.100 1.270 ;
        RECT  0.970 1.710 1.480 1.830 ;
        RECT  1.480 1.710 1.600 2.050 ;
        RECT  1.600 1.930 2.210 2.050 ;
        RECT  0.060 0.450 0.280 0.870 ;
        RECT  0.280 1.640 0.420 1.800 ;
        RECT  0.280 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.060 0.720 1.280 ;
        RECT  4.310 0.470 4.700 0.590 ;
        RECT  4.090 0.430 4.310 0.590 ;
        RECT  3.520 0.470 4.090 0.590 ;
        RECT  3.400 0.470 3.520 0.730 ;
        RECT  2.390 0.610 3.400 0.730 ;
        RECT  6.280 1.030 6.440 1.500 ;
        RECT  5.410 1.380 6.280 1.500 ;
        RECT  5.250 1.020 5.410 1.500 ;
        RECT  5.230 1.380 5.250 1.500 ;
        RECT  5.110 1.380 5.230 1.870 ;
        RECT  4.670 1.750 5.110 1.870 ;
        RECT  4.630 1.750 4.670 2.100 ;
        RECT  4.510 1.210 4.630 2.100 ;
        RECT  4.470 1.210 4.510 1.330 ;
        RECT  4.350 0.710 4.470 1.330 ;
        RECT  7.600 1.080 7.720 1.240 ;
        RECT  7.480 0.470 7.600 1.480 ;
        RECT  7.280 0.470 7.480 0.590 ;
        RECT  7.430 1.360 7.480 1.480 ;
        RECT  7.310 1.360 7.430 1.650 ;
        RECT  6.860 1.490 7.310 1.650 ;
        RECT  7.060 0.420 7.280 0.590 ;
        RECT  5.660 0.470 7.060 0.590 ;
        RECT  5.540 0.470 5.660 0.830 ;
        RECT  4.880 0.710 5.540 0.830 ;
        RECT  4.880 1.460 4.990 1.620 ;
        RECT  4.760 0.710 4.880 1.620 ;
        RECT  8.910 1.080 9.280 1.240 ;
        RECT  8.790 1.080 8.910 2.050 ;
        RECT  7.380 1.930 8.790 2.050 ;
        RECT  7.260 1.770 7.380 2.050 ;
        RECT  6.740 1.770 7.260 1.890 ;
        RECT  6.740 0.710 6.770 1.270 ;
        RECT  6.620 0.710 6.740 1.890 ;
        RECT  5.780 0.710 6.620 0.870 ;
        RECT  5.390 1.620 6.620 1.780 ;
        RECT  4.590 0.710 4.760 0.850 ;
        RECT  4.210 0.710 4.350 0.850 ;
        RECT  2.230 0.610 2.390 0.960 ;
        RECT  2.900 1.880 3.110 2.100 ;
        RECT  3.410 1.500 3.640 1.660 ;
        RECT  1.770 1.490 1.940 1.650 ;
        RECT  2.190 1.650 2.290 1.810 ;
        RECT  0.750 1.640 0.850 2.060 ;
        RECT  0.060 1.640 0.280 2.060 ;
        LAYER M1 ;
        RECT  9.160 1.650 9.335 2.030 ;
        RECT  9.160 0.490 9.335 0.870 ;
        RECT  8.585 0.490 8.640 0.870 ;
        RECT  7.720 0.490 7.735 0.870 ;
        RECT  7.570 1.600 7.735 1.760 ;
    END
END DFNCSND4

MACRO DFND1
    CLASS CORE ;
    FOREIGN DFND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.480 1.960 5.510 2.100 ;
        RECT  5.510 0.420 5.670 2.100 ;
        RECT  5.670 1.960 5.700 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.960 4.710 2.100 ;
        RECT  4.710 1.390 4.870 2.100 ;
        RECT  4.870 1.390 4.890 1.515 ;
        RECT  4.720 0.710 4.890 0.870 ;
        RECT  4.870 1.960 4.900 2.100 ;
        RECT  4.890 0.710 5.030 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.030 2.820 ;
        RECT  1.030 2.030 1.250 2.820 ;
        RECT  1.250 2.220 2.320 2.820 ;
        RECT  2.320 2.030 2.540 2.820 ;
        RECT  2.540 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.470 3.720 1.050 ;
        RECT  3.720 0.470 3.810 1.810 ;
        RECT  3.810 0.950 3.840 1.810 ;
        RECT  3.810 0.470 5.240 0.590 ;
        RECT  5.240 0.470 5.380 1.290 ;
        RECT  5.380 1.050 5.390 1.290 ;
        RECT  4.350 1.610 4.470 2.090 ;
        RECT  4.100 0.710 4.470 0.850 ;
        RECT  4.470 0.710 4.510 2.090 ;
        RECT  4.510 0.710 4.590 1.730 ;
        RECT  4.590 0.710 4.600 1.270 ;
        RECT  4.600 1.050 4.770 1.270 ;
        RECT  3.290 1.930 4.110 2.050 ;
        RECT  4.110 1.290 4.230 2.050 ;
        RECT  4.230 1.290 4.350 1.450 ;
        RECT  1.370 0.470 1.900 0.590 ;
        RECT  1.900 0.430 2.120 0.590 ;
        RECT  2.120 0.470 2.970 0.590 ;
        RECT  2.970 0.430 3.190 0.590 ;
        RECT  3.190 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.460 1.290 ;
        RECT  3.460 0.470 3.530 1.540 ;
        RECT  3.530 1.170 3.600 1.540 ;
        RECT  2.700 1.750 2.860 1.910 ;
        RECT  2.430 0.760 2.860 0.920 ;
        RECT  2.860 0.760 2.980 1.910 ;
        RECT  1.700 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  2.070 1.510 2.590 1.630 ;
        RECT  2.590 1.060 2.740 1.630 ;
        RECT  0.760 0.430 0.890 0.850 ;
        RECT  0.890 0.430 0.950 1.880 ;
        RECT  0.950 0.430 0.980 1.650 ;
        RECT  0.980 0.730 1.050 1.650 ;
        RECT  1.050 1.530 1.410 1.650 ;
        RECT  1.410 1.530 1.530 2.050 ;
        RECT  1.530 1.930 1.920 2.050 ;
        RECT  1.920 1.930 2.160 2.090 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.290 1.640 0.420 1.760 ;
        RECT  0.290 0.760 0.420 0.880 ;
        RECT  0.420 0.760 0.540 1.760 ;
        RECT  0.540 1.080 0.760 1.240 ;
        RECT  3.960 0.710 4.100 1.160 ;
        RECT  3.130 0.710 3.290 2.050 ;
        RECT  1.210 0.470 1.370 1.410 ;
        RECT  2.270 0.760 2.430 1.320 ;
        RECT  1.720 1.640 1.950 1.800 ;
        RECT  0.790 1.380 0.890 1.880 ;
        RECT  0.070 1.640 0.290 2.060 ;
        RECT  3.580 1.660 3.720 1.810 ;
    END
END DFND1

MACRO DFND2
    CLASS CORE ;
    FOREIGN DFND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.060 1.940 6.090 2.100 ;
        RECT  6.090 1.390 6.170 2.100 ;
        RECT  6.090 0.420 6.170 0.900 ;
        RECT  6.170 0.420 6.250 2.100 ;
        RECT  6.250 1.940 6.280 2.100 ;
        RECT  6.250 0.780 6.310 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.350 1.940 5.380 2.100 ;
        RECT  5.380 1.390 5.530 2.100 ;
        RECT  5.330 0.710 5.530 0.870 ;
        RECT  5.530 0.710 5.540 2.100 ;
        RECT  5.540 1.940 5.570 2.100 ;
        RECT  5.540 0.710 5.670 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 4.210 0.300 ;
        RECT  4.210 -0.300 4.430 0.340 ;
        RECT  4.430 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.410 2.820 ;
        RECT  2.410 2.030 2.630 2.820 ;
        RECT  2.630 2.220 4.210 2.820 ;
        RECT  4.210 2.180 4.430 2.820 ;
        RECT  4.430 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.380 1.930 4.250 2.050 ;
        RECT  4.250 1.390 4.370 2.050 ;
        RECT  4.370 1.390 4.570 1.510 ;
        RECT  4.570 1.030 4.730 1.510 ;
        RECT  0.070 0.720 0.420 0.880 ;
        RECT  0.420 0.510 0.540 1.950 ;
        RECT  0.540 0.510 0.750 0.630 ;
        RECT  0.750 0.470 0.845 0.630 ;
        RECT  0.540 1.115 0.850 1.275 ;
        RECT  0.845 0.470 1.900 0.590 ;
        RECT  1.900 0.430 2.120 0.590 ;
        RECT  2.120 0.470 3.515 0.590 ;
        RECT  3.515 0.470 3.635 1.540 ;
        RECT  3.635 1.320 3.680 1.540 ;
        RECT  2.790 1.750 2.905 1.910 ;
        RECT  2.410 0.760 2.905 0.920 ;
        RECT  2.905 0.760 3.030 1.910 ;
        RECT  1.700 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.790 ;
        RECT  2.070 1.510 2.590 1.630 ;
        RECT  2.590 1.050 2.750 1.630 ;
        RECT  0.980 1.640 1.190 1.800 ;
        RECT  0.740 0.750 1.190 0.910 ;
        RECT  1.190 0.750 1.350 1.800 ;
        RECT  1.350 1.640 1.370 1.800 ;
        RECT  1.370 1.640 1.490 2.050 ;
        RECT  1.490 1.910 2.240 2.050 ;
        RECT  5.015 1.080 5.410 1.240 ;
        RECT  5.010 0.710 5.015 1.240 ;
        RECT  4.850 0.710 5.010 1.750 ;
        RECT  4.310 0.710 4.850 0.870 ;
        RECT  4.845 1.630 4.850 1.750 ;
        RECT  4.625 1.630 4.845 2.050 ;
        RECT  5.950 1.080 6.050 1.240 ;
        RECT  5.830 0.470 5.950 1.240 ;
        RECT  4.010 0.470 5.830 0.590 ;
        RECT  3.860 0.470 4.010 1.810 ;
        RECT  4.170 0.710 4.310 1.270 ;
        RECT  3.220 0.710 3.380 2.050 ;
        RECT  0.070 1.790 0.420 1.950 ;
        RECT  2.250 0.760 2.410 1.320 ;
        RECT  1.720 1.635 1.950 1.790 ;
        RECT  0.760 1.640 0.980 2.060 ;
        RECT  3.650 1.660 3.860 1.810 ;
    END
END DFND2

MACRO DFND4
    CLASS CORE ;
    FOREIGN DFND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.310 1.650 7.630 2.030 ;
        RECT  7.310 0.510 7.630 0.890 ;
        RECT  7.630 0.510 8.050 2.030 ;
        RECT  8.050 1.650 8.220 2.030 ;
        RECT  8.050 0.510 8.220 0.890 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.930 1.650 6.350 2.030 ;
        RECT  5.910 0.760 6.350 0.920 ;
        RECT  6.350 0.760 6.770 2.030 ;
        RECT  6.770 1.650 6.840 2.030 ;
        RECT  6.770 0.760 6.860 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.030 0.300 ;
        RECT  1.030 -0.300 1.250 0.340 ;
        RECT  1.250 -0.300 2.430 0.300 ;
        RECT  2.430 -0.300 2.650 0.340 ;
        RECT  2.650 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.430 2.820 ;
        RECT  2.430 2.030 2.650 2.820 ;
        RECT  2.650 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 0.430 2.140 0.590 ;
        RECT  2.140 0.470 3.620 0.590 ;
        RECT  3.620 0.470 3.760 1.540 ;
        RECT  3.760 1.320 3.810 1.540 ;
        RECT  2.810 1.750 2.940 1.910 ;
        RECT  2.500 0.710 2.940 0.870 ;
        RECT  2.940 0.710 3.060 1.910 ;
        RECT  1.720 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.775 ;
        RECT  2.070 1.510 2.660 1.630 ;
        RECT  2.660 1.030 2.820 1.630 ;
        RECT  0.980 1.890 1.210 2.050 ;
        RECT  0.740 0.710 1.210 0.870 ;
        RECT  1.210 0.710 1.370 2.050 ;
        RECT  1.370 1.895 2.240 2.050 ;
        RECT  0.540 0.470 1.920 0.590 ;
        RECT  0.540 1.105 0.850 1.275 ;
        RECT  0.420 0.470 0.540 1.760 ;
        RECT  0.290 0.470 0.420 0.850 ;
        RECT  0.290 1.640 0.420 1.760 ;
        RECT  0.070 0.430 0.290 0.850 ;
        RECT  5.270 1.030 5.430 1.480 ;
        RECT  5.085 1.360 5.270 1.480 ;
        RECT  4.965 1.360 5.085 2.010 ;
        RECT  3.400 1.890 4.965 2.010 ;
        RECT  5.700 1.080 6.040 1.240 ;
        RECT  5.580 0.710 5.700 1.750 ;
        RECT  5.045 0.710 5.580 0.870 ;
        RECT  5.430 1.600 5.580 1.750 ;
        RECT  5.270 1.600 5.430 2.100 ;
        RECT  4.925 0.710 5.045 1.240 ;
        RECT  7.190 1.080 7.400 1.240 ;
        RECT  7.070 0.470 7.190 1.240 ;
        RECT  4.780 0.470 7.070 0.590 ;
        RECT  4.120 1.610 4.830 1.770 ;
        RECT  4.620 0.470 4.780 0.840 ;
        RECT  4.120 0.650 4.620 0.840 ;
        RECT  3.980 0.650 4.120 1.770 ;
        RECT  3.900 0.650 3.980 0.840 ;
        RECT  4.245 1.080 4.925 1.240 ;
        RECT  3.930 1.540 3.980 1.770 ;
        RECT  3.240 0.710 3.400 2.010 ;
        RECT  0.070 1.640 0.290 2.060 ;
        RECT  2.340 0.710 2.500 1.320 ;
        RECT  1.720 1.635 1.950 1.775 ;
        RECT  0.760 1.630 0.980 2.050 ;
        LAYER M1 ;
        RECT  5.910 0.760 6.135 0.920 ;
        RECT  5.930 1.650 6.135 2.030 ;
        RECT  7.310 1.650 7.415 2.030 ;
        RECT  7.310 0.510 7.415 0.890 ;
    END
END DFND4

MACRO DFNSND1
    CLASS CORE ;
    FOREIGN DFNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 1.940 6.470 2.100 ;
        RECT  6.470 1.390 6.510 2.100 ;
        RECT  6.470 0.420 6.510 0.900 ;
        RECT  6.510 0.420 6.650 2.100 ;
        RECT  6.650 1.940 6.660 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.750 1.940 5.780 2.100 ;
        RECT  5.780 1.390 5.850 2.100 ;
        RECT  5.750 0.710 5.850 0.870 ;
        RECT  5.850 0.710 5.940 2.100 ;
        RECT  5.940 1.940 5.970 2.100 ;
        RECT  5.940 0.710 5.990 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.080 1.790 1.240 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 0.990 0.300 ;
        RECT  0.990 -0.300 1.210 0.480 ;
        RECT  1.210 -0.300 2.410 0.300 ;
        RECT  2.410 -0.300 2.630 0.340 ;
        RECT  2.630 -0.300 4.990 0.300 ;
        RECT  4.990 -0.300 5.210 0.340 ;
        RECT  5.210 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 0.990 2.820 ;
        RECT  0.990 1.990 1.210 2.820 ;
        RECT  1.210 2.220 2.270 2.820 ;
        RECT  2.270 2.170 2.490 2.820 ;
        RECT  2.490 2.220 3.070 2.820 ;
        RECT  3.070 2.060 3.290 2.820 ;
        RECT  3.290 2.220 4.310 2.820 ;
        RECT  4.310 1.980 4.530 2.820 ;
        RECT  4.530 2.220 5.000 2.820 ;
        RECT  5.000 2.180 5.220 2.820 ;
        RECT  5.220 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.530 0.470 4.000 0.590 ;
        RECT  4.000 0.430 4.240 0.590 ;
        RECT  0.730 0.680 0.870 0.840 ;
        RECT  0.870 0.680 0.990 1.800 ;
        RECT  0.990 1.010 1.180 1.230 ;
        RECT  0.990 1.680 1.360 1.800 ;
        RECT  1.360 1.680 1.480 2.050 ;
        RECT  1.480 1.930 1.890 2.050 ;
        RECT  1.890 1.930 2.110 2.090 ;
        RECT  2.110 1.930 2.280 2.050 ;
        RECT  2.280 1.820 2.400 2.050 ;
        RECT  2.400 1.820 3.410 1.940 ;
        RECT  3.410 1.820 3.530 2.100 ;
        RECT  3.530 1.960 3.650 2.100 ;
        RECT  2.360 1.580 3.090 1.700 ;
        RECT  3.090 0.710 3.250 1.700 ;
        RECT  3.250 1.560 3.550 1.700 ;
        RECT  1.700 0.710 1.910 0.850 ;
        RECT  1.910 0.710 2.030 1.810 ;
        RECT  2.030 1.030 2.520 1.150 ;
        RECT  2.520 1.030 2.680 1.340 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.080 0.750 1.240 ;
        RECT  3.310 0.430 3.530 0.590 ;
        RECT  2.110 0.470 3.310 0.590 ;
        RECT  5.280 1.050 5.390 1.270 ;
        RECT  5.160 1.050 5.280 1.860 ;
        RECT  3.880 1.740 5.160 1.860 ;
        RECT  3.720 1.320 3.880 1.860 ;
        RECT  3.650 1.320 3.720 1.440 ;
        RECT  5.630 1.050 5.730 1.270 ;
        RECT  5.510 0.710 5.630 1.740 ;
        RECT  5.030 0.710 5.510 0.870 ;
        RECT  5.400 1.580 5.510 1.740 ;
        RECT  6.340 1.050 6.390 1.290 ;
        RECT  6.220 0.470 6.340 1.290 ;
        RECT  4.520 0.470 6.220 0.590 ;
        RECT  4.120 1.460 4.950 1.620 ;
        RECT  4.360 0.470 4.520 0.870 ;
        RECT  4.120 0.710 4.360 0.870 ;
        RECT  4.000 0.710 4.120 1.620 ;
        RECT  4.870 0.710 5.030 1.290 ;
        RECT  3.500 0.710 3.650 1.440 ;
        RECT  1.870 0.430 2.110 0.590 ;
        RECT  0.730 1.640 0.870 1.800 ;
        RECT  2.200 1.270 2.360 1.700 ;
        RECT  1.680 1.650 1.910 1.810 ;
        RECT  0.060 1.640 0.420 1.800 ;
        RECT  3.830 0.710 4.000 0.870 ;
    END
END DFNSND1

MACRO DFNSND2
    CLASS CORE ;
    FOREIGN DFNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.725 3.110 1.320 ;
        RECT  3.110 1.100 3.260 1.320 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.040 1.940 7.070 2.100 ;
        RECT  7.070 1.390 7.130 2.100 ;
        RECT  7.070 0.420 7.130 0.900 ;
        RECT  7.130 0.420 7.230 2.100 ;
        RECT  7.230 1.940 7.260 2.100 ;
        RECT  7.230 0.780 7.270 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.940 6.380 2.100 ;
        RECT  6.380 1.390 6.490 2.100 ;
        RECT  6.330 0.710 6.490 0.870 ;
        RECT  6.490 0.710 6.540 2.100 ;
        RECT  6.540 1.940 6.570 2.100 ;
        RECT  6.540 0.710 6.630 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.925 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.110 0.300 ;
        RECT  1.110 -0.300 1.330 0.480 ;
        RECT  1.330 -0.300 2.550 0.300 ;
        RECT  2.550 -0.300 2.770 0.340 ;
        RECT  2.770 -0.300 5.140 0.300 ;
        RECT  5.140 -0.300 5.360 0.340 ;
        RECT  5.360 -0.300 5.960 0.300 ;
        RECT  5.960 -0.300 6.180 0.340 ;
        RECT  6.180 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.100 2.820 ;
        RECT  1.100 1.990 1.320 2.820 ;
        RECT  1.320 2.220 2.420 2.820 ;
        RECT  2.420 2.170 2.640 2.820 ;
        RECT  2.640 2.220 3.220 2.820 ;
        RECT  3.220 2.060 3.440 2.820 ;
        RECT  3.440 2.220 4.460 2.820 ;
        RECT  4.460 1.980 4.680 2.820 ;
        RECT  4.680 2.220 5.960 2.820 ;
        RECT  5.960 2.180 6.180 2.820 ;
        RECT  6.180 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.750 1.240 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  2.650 1.010 2.810 1.340 ;
        RECT  2.180 1.010 2.650 1.130 ;
        RECT  2.060 0.710 2.180 1.785 ;
        RECT  1.820 0.710 2.060 0.870 ;
        RECT  3.500 1.560 3.700 1.700 ;
        RECT  3.380 0.710 3.500 1.700 ;
        RECT  3.290 0.710 3.380 0.930 ;
        RECT  2.490 1.520 3.380 1.700 ;
        RECT  3.680 1.960 3.800 2.100 ;
        RECT  3.560 1.820 3.680 2.100 ;
        RECT  2.550 1.820 3.560 1.940 ;
        RECT  2.430 1.820 2.550 2.025 ;
        RECT  2.260 1.905 2.430 2.025 ;
        RECT  2.040 1.905 2.260 2.060 ;
        RECT  1.590 1.905 2.040 2.025 ;
        RECT  1.470 1.680 1.590 2.025 ;
        RECT  0.990 1.020 1.510 1.180 ;
        RECT  0.990 1.680 1.470 1.800 ;
        RECT  0.970 0.710 0.990 1.800 ;
        RECT  0.870 0.710 0.970 2.060 ;
        RECT  0.730 0.710 0.870 0.870 ;
        RECT  4.170 0.430 4.390 0.590 ;
        RECT  2.265 0.470 4.170 0.590 ;
        RECT  5.460 1.050 5.540 1.270 ;
        RECT  5.340 1.050 5.460 1.860 ;
        RECT  4.030 1.740 5.340 1.860 ;
        RECT  3.870 1.320 4.030 1.860 ;
        RECT  3.850 1.320 3.870 1.440 ;
        RECT  5.780 1.080 6.370 1.240 ;
        RECT  5.740 0.710 5.780 1.700 ;
        RECT  5.660 0.710 5.740 2.080 ;
        RECT  5.180 0.710 5.660 0.870 ;
        RECT  5.580 1.580 5.660 2.080 ;
        RECT  6.950 1.050 7.010 1.270 ;
        RECT  6.830 0.470 6.950 1.270 ;
        RECT  4.670 0.470 6.830 0.590 ;
        RECT  4.670 1.460 5.100 1.620 ;
        RECT  4.510 0.470 4.670 1.620 ;
        RECT  4.030 0.710 4.510 0.870 ;
        RECT  5.020 0.710 5.180 1.290 ;
        RECT  3.690 0.710 3.850 1.440 ;
        RECT  2.025 0.430 2.265 0.590 ;
        RECT  0.750 1.640 0.870 2.060 ;
        RECT  2.330 1.250 2.490 1.700 ;
        RECT  1.810 1.635 2.060 1.785 ;
        RECT  0.060 1.640 0.420 1.800 ;
        RECT  4.200 1.460 4.510 1.620 ;
    END
END DFNSND2

MACRO DFNSND4
    CLASS CORE ;
    FOREIGN DFNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.725 3.110 1.320 ;
        RECT  3.110 1.100 3.270 1.320 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.810 1.650 8.270 2.030 ;
        RECT  7.810 0.490 8.270 0.870 ;
        RECT  8.270 0.490 8.690 2.030 ;
        RECT  8.690 1.650 8.750 2.030 ;
        RECT  8.690 0.490 8.750 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.370 1.650 6.670 2.030 ;
        RECT  6.350 0.760 6.670 0.920 ;
        RECT  6.670 0.760 7.090 2.030 ;
        RECT  7.090 1.650 7.310 2.030 ;
        RECT  7.090 0.760 7.330 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.920 1.270 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.110 0.300 ;
        RECT  1.110 -0.300 1.330 0.480 ;
        RECT  1.330 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 5.120 0.300 ;
        RECT  5.120 -0.300 5.340 0.340 ;
        RECT  5.340 -0.300 5.970 0.300 ;
        RECT  5.970 -0.300 6.190 0.340 ;
        RECT  6.190 -0.300 8.930 0.300 ;
        RECT  8.930 -0.300 9.150 0.340 ;
        RECT  9.150 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.100 2.820 ;
        RECT  1.100 1.990 1.320 2.820 ;
        RECT  1.320 2.220 2.400 2.820 ;
        RECT  2.400 2.180 2.620 2.820 ;
        RECT  2.620 2.220 3.200 2.820 ;
        RECT  3.200 2.060 3.420 2.820 ;
        RECT  3.420 2.220 4.440 2.820 ;
        RECT  4.440 1.980 4.660 2.820 ;
        RECT  4.660 2.220 5.970 2.820 ;
        RECT  5.970 2.170 6.190 2.820 ;
        RECT  6.190 2.220 8.930 2.820 ;
        RECT  8.930 2.170 9.155 2.820 ;
        RECT  9.155 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.750 1.240 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.280 0.710 0.420 0.870 ;
        RECT  0.280 1.640 0.420 1.800 ;
        RECT  0.060 0.450 0.280 0.870 ;
        RECT  2.630 1.010 2.790 1.340 ;
        RECT  2.160 1.010 2.630 1.130 ;
        RECT  2.040 0.710 2.160 1.795 ;
        RECT  1.800 0.710 2.040 0.870 ;
        RECT  3.510 1.560 3.680 1.700 ;
        RECT  3.390 0.740 3.510 1.700 ;
        RECT  3.240 0.740 3.390 0.900 ;
        RECT  2.470 1.550 3.390 1.700 ;
        RECT  3.660 1.960 3.780 2.100 ;
        RECT  3.540 1.820 3.660 2.100 ;
        RECT  2.530 1.820 3.540 1.940 ;
        RECT  2.410 1.820 2.530 2.050 ;
        RECT  2.240 1.930 2.410 2.050 ;
        RECT  2.020 1.930 2.240 2.070 ;
        RECT  1.570 1.930 2.020 2.050 ;
        RECT  1.450 1.680 1.570 2.050 ;
        RECT  0.990 0.935 1.500 1.110 ;
        RECT  0.990 1.680 1.450 1.800 ;
        RECT  0.970 0.710 0.990 1.800 ;
        RECT  0.870 0.450 0.970 2.060 ;
        RECT  0.750 0.450 0.870 0.870 ;
        RECT  4.150 0.430 4.370 0.590 ;
        RECT  2.245 0.470 4.150 0.590 ;
        RECT  5.440 1.050 5.520 1.270 ;
        RECT  5.320 1.050 5.440 1.860 ;
        RECT  4.010 1.740 5.320 1.860 ;
        RECT  3.850 1.320 4.010 1.860 ;
        RECT  3.830 1.320 3.850 1.440 ;
        RECT  5.760 1.080 6.410 1.240 ;
        RECT  5.720 0.710 5.760 1.510 ;
        RECT  5.720 1.960 5.750 2.100 ;
        RECT  5.640 0.710 5.720 2.100 ;
        RECT  5.160 0.710 5.640 0.870 ;
        RECT  5.560 1.390 5.640 2.100 ;
        RECT  5.530 1.960 5.560 2.100 ;
        RECT  7.635 1.080 7.920 1.240 ;
        RECT  7.515 0.470 7.635 1.240 ;
        RECT  4.650 0.470 7.515 0.590 ;
        RECT  4.650 1.460 5.080 1.620 ;
        RECT  4.490 0.470 4.650 1.620 ;
        RECT  4.010 0.710 4.490 0.870 ;
        RECT  5.000 0.710 5.160 1.290 ;
        RECT  3.670 0.710 3.830 1.440 ;
        RECT  2.005 0.430 2.245 0.590 ;
        RECT  0.750 1.640 0.870 2.060 ;
        RECT  2.310 1.250 2.470 1.700 ;
        RECT  1.790 1.635 2.040 1.795 ;
        RECT  4.180 1.480 4.490 1.620 ;
        RECT  0.060 1.640 0.280 2.060 ;
        LAYER M1 ;
        RECT  7.810 0.490 8.055 0.870 ;
        RECT  7.305 1.650 7.310 2.030 ;
        RECT  7.305 0.760 7.330 0.920 ;
        RECT  6.370 1.650 6.455 2.030 ;
        RECT  6.350 0.760 6.455 0.920 ;
        RECT  7.810 1.650 8.055 2.030 ;
    END
END DFNSND4

MACRO DFQD1
    CLASS CORE ;
    FOREIGN DFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.680 1.960 4.710 2.100 ;
        RECT  4.710 1.390 4.870 2.100 ;
        RECT  4.870 1.390 4.890 1.515 ;
        RECT  4.770 0.420 4.890 0.900 ;
        RECT  4.870 1.960 4.900 2.100 ;
        RECT  4.890 0.420 4.930 1.515 ;
        RECT  4.930 0.780 5.030 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.020 2.820 ;
        RECT  1.020 2.030 1.240 2.820 ;
        RECT  1.240 2.220 2.320 2.820 ;
        RECT  2.320 2.030 2.540 2.820 ;
        RECT  2.540 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.190 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.460 1.290 ;
        RECT  3.460 0.470 3.530 1.540 ;
        RECT  3.530 1.170 3.600 1.540 ;
        RECT  2.700 1.750 2.860 1.910 ;
        RECT  2.390 0.760 2.860 0.920 ;
        RECT  2.860 0.760 2.980 1.910 ;
        RECT  1.690 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  2.070 1.510 2.580 1.630 ;
        RECT  2.580 1.060 2.740 1.630 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.290 1.640 0.420 1.760 ;
        RECT  0.290 0.760 0.420 0.880 ;
        RECT  0.420 0.760 0.540 1.760 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  2.970 0.430 3.190 0.590 ;
        RECT  2.110 0.470 2.970 0.590 ;
        RECT  1.890 0.430 2.110 0.590 ;
        RECT  1.510 0.470 1.890 0.590 ;
        RECT  1.390 0.470 1.510 0.850 ;
        RECT  1.350 0.690 1.390 0.850 ;
        RECT  1.190 0.690 1.350 1.530 ;
        RECT  0.980 0.690 1.190 0.850 ;
        RECT  0.980 1.410 1.190 1.530 ;
        RECT  0.760 0.430 0.980 0.850 ;
        RECT  3.810 0.950 3.840 1.810 ;
        RECT  3.720 0.620 3.810 1.810 ;
        RECT  3.650 0.620 3.720 1.050 ;
        RECT  4.230 1.290 4.350 1.450 ;
        RECT  4.110 1.290 4.230 2.050 ;
        RECT  3.290 1.930 4.110 2.050 ;
        RECT  4.600 1.050 4.770 1.270 ;
        RECT  4.590 0.430 4.600 1.270 ;
        RECT  4.510 0.430 4.590 1.730 ;
        RECT  4.470 0.430 4.510 2.090 ;
        RECT  4.380 0.430 4.470 0.850 ;
        RECT  4.350 1.610 4.470 2.090 ;
        RECT  4.100 0.730 4.380 0.850 ;
        RECT  3.130 0.710 3.290 2.050 ;
        RECT  3.580 1.660 3.720 1.810 ;
        RECT  0.760 1.410 0.980 1.830 ;
        RECT  2.230 0.760 2.390 1.320 ;
        RECT  1.700 1.640 1.950 1.800 ;
        RECT  0.070 1.640 0.290 2.060 ;
        RECT  3.960 0.730 4.100 1.160 ;
    END
END DFQD1

MACRO DFQD2
    CLASS CORE ;
    FOREIGN DFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.110 1.950 5.140 2.090 ;
        RECT  5.140 1.380 5.300 2.090 ;
        RECT  5.140 0.420 5.300 0.920 ;
        RECT  5.300 1.950 5.330 2.090 ;
        RECT  5.300 1.380 5.530 1.515 ;
        RECT  5.300 0.800 5.530 0.920 ;
        RECT  5.530 0.800 5.670 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.340 ;
        RECT  0.580 -0.300 2.310 0.300 ;
        RECT  2.310 -0.300 2.530 0.340 ;
        RECT  2.530 -0.300 3.990 0.300 ;
        RECT  3.990 -0.300 4.210 0.360 ;
        RECT  4.210 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.020 2.820 ;
        RECT  1.020 2.030 1.240 2.820 ;
        RECT  1.240 2.220 2.270 2.820 ;
        RECT  2.270 2.030 2.490 2.820 ;
        RECT  2.490 2.220 4.000 2.820 ;
        RECT  4.000 2.180 4.220 2.820 ;
        RECT  4.220 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  0.420 0.710 0.540 1.795 ;
        RECT  0.070 0.710 0.420 0.870 ;
        RECT  2.550 1.060 2.710 1.630 ;
        RECT  2.070 1.510 2.550 1.630 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  1.680 0.710 1.950 0.870 ;
        RECT  2.830 0.760 2.950 1.910 ;
        RECT  2.390 0.760 2.830 0.920 ;
        RECT  2.650 1.750 2.830 1.910 ;
        RECT  3.480 0.470 3.600 1.560 ;
        RECT  3.120 0.470 3.480 0.590 ;
        RECT  3.460 1.290 3.480 1.560 ;
        RECT  2.900 0.450 3.120 0.590 ;
        RECT  2.120 0.470 2.900 0.590 ;
        RECT  1.900 0.430 2.120 0.590 ;
        RECT  1.550 0.470 1.900 0.590 ;
        RECT  1.390 0.470 1.550 0.850 ;
        RECT  1.350 0.690 1.390 0.850 ;
        RECT  1.190 0.690 1.350 1.530 ;
        RECT  0.980 0.690 1.190 0.850 ;
        RECT  0.980 1.410 1.190 1.530 ;
        RECT  0.760 0.430 0.980 0.850 ;
        RECT  4.270 1.030 4.430 1.510 ;
        RECT  4.140 1.390 4.270 1.510 ;
        RECT  4.020 1.390 4.140 2.050 ;
        RECT  3.280 1.930 4.020 2.050 ;
        RECT  4.790 1.080 5.220 1.240 ;
        RECT  4.670 0.710 4.790 1.750 ;
        RECT  4.050 0.710 4.670 0.870 ;
        RECT  4.610 1.630 4.670 1.750 ;
        RECT  4.390 1.630 4.610 2.050 ;
        RECT  3.910 0.710 4.050 1.270 ;
        RECT  3.120 0.710 3.280 2.050 ;
        RECT  0.760 1.410 0.980 1.830 ;
        RECT  2.230 0.760 2.390 1.320 ;
        RECT  1.700 1.640 1.950 1.800 ;
        RECT  0.070 1.635 0.420 1.795 ;
    END
END DFQD2

MACRO DFQD4
    CLASS CORE ;
    FOREIGN DFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.010 1.650 5.390 2.030 ;
        RECT  5.010 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.950 2.030 ;
        RECT  5.810 0.490 5.950 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.310 0.300 ;
        RECT  2.310 -0.300 2.530 0.340 ;
        RECT  2.530 -0.300 3.910 0.300 ;
        RECT  3.910 -0.300 4.130 0.340 ;
        RECT  4.130 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.020 2.820 ;
        RECT  1.020 2.030 1.240 2.820 ;
        RECT  1.240 2.220 2.270 2.820 ;
        RECT  2.270 2.030 2.490 2.820 ;
        RECT  2.490 2.220 3.910 2.820 ;
        RECT  3.910 2.180 4.130 2.820 ;
        RECT  4.130 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.850 1.240 ;
        RECT  0.420 0.760 0.540 1.760 ;
        RECT  0.290 0.760 0.420 0.880 ;
        RECT  0.290 1.640 0.420 1.760 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  2.550 1.060 2.710 1.630 ;
        RECT  2.070 1.510 2.550 1.630 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  1.700 0.710 1.950 0.870 ;
        RECT  2.830 0.760 2.950 1.910 ;
        RECT  2.390 0.760 2.830 0.920 ;
        RECT  2.650 1.750 2.830 1.910 ;
        RECT  3.450 0.470 3.610 1.560 ;
        RECT  3.120 0.470 3.450 0.590 ;
        RECT  2.900 0.450 3.120 0.590 ;
        RECT  2.120 0.470 2.900 0.590 ;
        RECT  1.900 0.430 2.120 0.590 ;
        RECT  1.510 0.470 1.900 0.590 ;
        RECT  1.390 0.470 1.510 0.850 ;
        RECT  1.350 0.690 1.390 0.850 ;
        RECT  1.190 0.690 1.350 1.530 ;
        RECT  0.980 0.690 1.190 0.850 ;
        RECT  0.980 1.410 1.190 1.530 ;
        RECT  0.760 0.430 0.980 0.850 ;
        RECT  4.340 1.030 4.500 1.510 ;
        RECT  4.140 1.390 4.340 1.510 ;
        RECT  4.020 1.390 4.140 2.050 ;
        RECT  3.280 1.930 4.020 2.050 ;
        RECT  4.790 1.080 5.120 1.240 ;
        RECT  4.670 0.750 4.790 1.750 ;
        RECT  4.530 0.750 4.670 0.870 ;
        RECT  4.530 1.630 4.670 1.750 ;
        RECT  4.310 0.450 4.530 0.870 ;
        RECT  4.310 1.630 4.530 2.050 ;
        RECT  3.950 0.750 4.310 0.870 ;
        RECT  3.120 0.710 3.280 2.050 ;
        RECT  0.760 1.410 0.980 1.830 ;
        RECT  2.230 0.760 2.390 1.320 ;
        RECT  1.700 1.640 1.950 1.800 ;
        RECT  0.070 1.640 0.290 2.060 ;
        RECT  3.790 0.750 3.950 1.270 ;
        LAYER M1 ;
        RECT  5.010 1.650 5.175 2.030 ;
        RECT  5.010 0.490 5.175 0.870 ;
    END
END DFQD4

MACRO DFSND1
    CLASS CORE ;
    FOREIGN DFSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 1.940 6.470 2.100 ;
        RECT  6.470 1.390 6.510 2.100 ;
        RECT  6.470 0.420 6.510 0.900 ;
        RECT  6.510 0.420 6.630 2.100 ;
        RECT  6.630 1.940 6.660 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.750 1.940 5.780 2.100 ;
        RECT  5.780 1.390 5.850 2.100 ;
        RECT  5.750 0.710 5.850 0.870 ;
        RECT  5.850 0.710 5.940 2.100 ;
        RECT  5.940 1.940 5.970 2.100 ;
        RECT  5.940 0.710 5.990 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.570 1.050 1.690 1.270 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 0.990 0.300 ;
        RECT  0.990 -0.300 1.210 0.480 ;
        RECT  1.210 -0.300 2.420 0.300 ;
        RECT  2.420 -0.300 2.640 0.340 ;
        RECT  2.640 -0.300 5.000 0.300 ;
        RECT  5.000 -0.300 5.220 0.340 ;
        RECT  5.220 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 0.990 2.820 ;
        RECT  0.990 1.990 1.210 2.820 ;
        RECT  1.210 2.220 2.280 2.820 ;
        RECT  2.280 2.170 2.500 2.820 ;
        RECT  2.500 2.220 3.080 2.820 ;
        RECT  3.080 2.060 3.300 2.820 ;
        RECT  3.300 2.220 4.320 2.820 ;
        RECT  4.320 1.980 4.540 2.820 ;
        RECT  4.540 2.220 5.010 2.820 ;
        RECT  5.010 2.180 5.230 2.820 ;
        RECT  5.230 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.730 0.710 0.870 0.870 ;
        RECT  0.870 0.710 0.990 1.800 ;
        RECT  0.990 1.240 1.380 1.400 ;
        RECT  0.990 0.710 1.410 0.830 ;
        RECT  1.410 0.470 1.530 0.830 ;
        RECT  1.530 0.470 3.320 0.590 ;
        RECT  3.320 0.430 3.540 0.590 ;
        RECT  3.540 0.470 4.010 0.590 ;
        RECT  4.010 0.430 4.250 0.590 ;
        RECT  2.120 1.920 2.290 2.040 ;
        RECT  2.290 1.820 2.410 2.040 ;
        RECT  2.410 1.820 3.420 1.940 ;
        RECT  3.420 1.820 3.540 2.100 ;
        RECT  3.540 1.960 3.660 2.100 ;
        RECT  2.360 1.560 3.100 1.700 ;
        RECT  3.100 0.710 3.260 1.700 ;
        RECT  3.260 1.560 3.560 1.700 ;
        RECT  1.720 0.710 1.950 0.870 ;
        RECT  1.950 0.710 2.070 1.800 ;
        RECT  2.070 0.960 2.560 1.080 ;
        RECT  2.560 0.960 2.720 1.340 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.080 0.750 1.240 ;
        RECT  5.320 1.050 5.390 1.270 ;
        RECT  5.200 1.050 5.320 1.860 ;
        RECT  3.890 1.740 5.200 1.860 ;
        RECT  3.730 1.320 3.890 1.860 ;
        RECT  3.660 1.320 3.730 1.440 ;
        RECT  5.630 1.050 5.730 1.270 ;
        RECT  5.600 0.710 5.630 1.620 ;
        RECT  5.510 0.710 5.600 2.000 ;
        RECT  5.040 0.710 5.510 0.870 ;
        RECT  5.440 1.500 5.510 2.000 ;
        RECT  6.340 1.050 6.390 1.290 ;
        RECT  6.220 0.470 6.340 1.290 ;
        RECT  4.530 0.470 6.220 0.590 ;
        RECT  4.130 1.460 4.960 1.620 ;
        RECT  4.370 0.470 4.530 0.870 ;
        RECT  4.130 0.710 4.370 0.870 ;
        RECT  4.010 0.710 4.130 1.620 ;
        RECT  3.840 0.710 4.010 0.870 ;
        RECT  4.880 0.710 5.040 1.290 ;
        RECT  3.520 0.710 3.660 1.440 ;
        RECT  0.730 1.640 0.870 1.800 ;
        RECT  1.880 1.920 2.120 2.080 ;
        RECT  2.220 1.200 2.360 1.700 ;
        RECT  1.680 1.640 1.950 1.800 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFSND1

MACRO DFSND2
    CLASS CORE ;
    FOREIGN DFSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.725 3.110 1.320 ;
        RECT  3.110 1.100 3.270 1.320 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.020 1.940 7.050 2.100 ;
        RECT  7.050 1.390 7.130 2.100 ;
        RECT  7.050 0.420 7.130 0.900 ;
        RECT  7.130 0.420 7.210 2.100 ;
        RECT  7.210 1.940 7.240 2.100 ;
        RECT  7.210 0.780 7.270 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.310 1.940 6.340 2.100 ;
        RECT  6.340 1.390 6.490 2.100 ;
        RECT  6.290 0.710 6.490 0.870 ;
        RECT  6.490 0.710 6.500 2.100 ;
        RECT  6.500 1.940 6.530 2.100 ;
        RECT  6.500 0.710 6.630 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.860 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 1.110 0.300 ;
        RECT  1.110 -0.300 1.330 0.480 ;
        RECT  1.330 -0.300 2.540 0.300 ;
        RECT  2.540 -0.300 2.760 0.340 ;
        RECT  2.760 -0.300 5.120 0.300 ;
        RECT  5.120 -0.300 5.340 0.340 ;
        RECT  5.340 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.350 2.820 ;
        RECT  0.350 2.180 0.570 2.820 ;
        RECT  0.570 2.220 1.100 2.820 ;
        RECT  1.100 1.990 1.320 2.820 ;
        RECT  1.320 2.220 2.400 2.820 ;
        RECT  2.400 2.170 2.620 2.820 ;
        RECT  2.620 2.220 3.200 2.820 ;
        RECT  3.200 2.060 3.420 2.820 ;
        RECT  3.420 2.220 4.440 2.820 ;
        RECT  4.440 1.980 4.660 2.820 ;
        RECT  4.660 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.630 1.010 2.790 1.340 ;
        RECT  0.060 0.710 0.420 0.870 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.540 1.080 0.770 1.240 ;
        RECT  2.160 1.010 2.630 1.130 ;
        RECT  2.040 0.710 2.160 1.810 ;
        RECT  1.820 0.710 2.040 0.870 ;
        RECT  3.510 1.560 3.680 1.700 ;
        RECT  3.390 0.710 3.510 1.700 ;
        RECT  3.290 0.710 3.390 0.930 ;
        RECT  2.470 1.550 3.390 1.700 ;
        RECT  3.660 1.960 3.780 2.100 ;
        RECT  3.540 1.820 3.660 2.100 ;
        RECT  2.530 1.820 3.540 1.940 ;
        RECT  2.410 1.820 2.530 2.050 ;
        RECT  2.240 1.930 2.410 2.050 ;
        RECT  4.150 0.430 4.370 0.590 ;
        RECT  1.690 0.470 4.150 0.590 ;
        RECT  1.510 0.470 1.690 0.870 ;
        RECT  1.370 0.710 1.510 0.870 ;
        RECT  1.210 0.710 1.370 1.800 ;
        RECT  0.730 0.710 1.210 0.870 ;
        RECT  0.970 1.640 1.210 1.800 ;
        RECT  5.440 1.050 5.520 1.270 ;
        RECT  5.320 1.050 5.440 1.860 ;
        RECT  4.010 1.740 5.320 1.860 ;
        RECT  3.850 1.320 4.010 1.860 ;
        RECT  3.830 1.320 3.850 1.440 ;
        RECT  5.760 1.080 6.350 1.240 ;
        RECT  5.720 0.710 5.760 1.700 ;
        RECT  5.640 0.710 5.720 2.080 ;
        RECT  5.160 0.710 5.640 0.870 ;
        RECT  5.560 1.580 5.640 2.080 ;
        RECT  6.930 1.050 6.990 1.270 ;
        RECT  6.810 0.470 6.930 1.270 ;
        RECT  4.650 0.470 6.810 0.590 ;
        RECT  4.650 1.460 5.080 1.620 ;
        RECT  4.490 0.470 4.650 1.620 ;
        RECT  4.010 0.710 4.490 0.870 ;
        RECT  4.180 1.480 4.490 1.620 ;
        RECT  5.000 0.710 5.160 1.290 ;
        RECT  3.680 0.710 3.830 1.440 ;
        RECT  0.750 1.640 0.970 2.060 ;
        RECT  2.000 1.930 2.240 2.090 ;
        RECT  2.310 1.250 2.470 1.700 ;
        RECT  1.790 1.650 2.040 1.810 ;
        RECT  0.060 1.640 0.420 1.800 ;
    END
END DFSND2

MACRO DFSND4
    CLASS CORE ;
    FOREIGN DFSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.725 3.110 1.310 ;
        RECT  3.110 1.090 3.280 1.310 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.890 1.650 8.270 2.030 ;
        RECT  7.890 0.490 8.270 0.870 ;
        RECT  8.270 0.490 8.690 2.030 ;
        RECT  8.690 1.650 8.830 2.030 ;
        RECT  8.690 0.490 8.830 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.360 1.650 6.670 2.030 ;
        RECT  6.340 0.760 6.670 0.920 ;
        RECT  6.670 0.760 7.090 2.030 ;
        RECT  7.090 1.650 7.390 2.030 ;
        RECT  7.090 0.760 7.410 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.110 0.300 ;
        RECT  1.110 -0.300 1.330 0.480 ;
        RECT  1.330 -0.300 2.545 0.300 ;
        RECT  2.545 -0.300 2.765 0.350 ;
        RECT  2.765 -0.300 5.120 0.300 ;
        RECT  5.120 -0.300 5.345 0.350 ;
        RECT  5.345 -0.300 5.960 0.300 ;
        RECT  5.960 -0.300 6.180 0.340 ;
        RECT  6.180 -0.300 6.770 0.300 ;
        RECT  6.770 -0.300 6.990 0.340 ;
        RECT  6.990 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.100 2.820 ;
        RECT  1.100 1.990 1.320 2.820 ;
        RECT  1.320 2.220 2.410 2.820 ;
        RECT  2.410 2.180 2.630 2.820 ;
        RECT  2.630 2.220 3.210 2.820 ;
        RECT  3.210 2.060 3.430 2.820 ;
        RECT  3.430 2.220 4.450 2.820 ;
        RECT  4.450 1.980 4.670 2.820 ;
        RECT  4.670 2.220 5.960 2.820 ;
        RECT  5.960 2.170 6.180 2.820 ;
        RECT  6.180 2.220 6.770 2.820 ;
        RECT  6.770 2.180 6.990 2.820 ;
        RECT  6.990 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.765 1.240 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.280 0.710 0.420 0.870 ;
        RECT  0.280 1.640 0.420 1.800 ;
        RECT  0.060 0.450 0.280 0.870 ;
        RECT  2.640 1.010 2.800 1.340 ;
        RECT  2.170 1.010 2.640 1.130 ;
        RECT  2.050 0.710 2.170 1.810 ;
        RECT  1.810 0.710 2.050 0.870 ;
        RECT  3.520 1.560 3.690 1.700 ;
        RECT  3.400 0.710 3.520 1.700 ;
        RECT  3.280 0.710 3.400 0.930 ;
        RECT  2.480 1.550 3.400 1.700 ;
        RECT  3.670 1.960 3.790 2.100 ;
        RECT  3.550 1.820 3.670 2.100 ;
        RECT  2.540 1.820 3.550 1.940 ;
        RECT  2.420 1.820 2.540 2.050 ;
        RECT  2.250 1.930 2.420 2.050 ;
        RECT  4.160 0.430 4.380 0.590 ;
        RECT  1.630 0.470 4.160 0.590 ;
        RECT  1.505 0.470 1.630 0.870 ;
        RECT  1.005 0.710 1.505 0.870 ;
        RECT  1.005 1.240 1.430 1.400 ;
        RECT  0.980 0.710 1.005 1.800 ;
        RECT  0.970 0.450 0.980 1.800 ;
        RECT  0.885 0.450 0.970 2.060 ;
        RECT  0.760 0.450 0.885 0.870 ;
        RECT  5.450 1.050 5.530 1.270 ;
        RECT  5.330 1.050 5.450 1.860 ;
        RECT  4.020 1.740 5.330 1.860 ;
        RECT  3.860 1.320 4.020 1.860 ;
        RECT  3.840 1.320 3.860 1.440 ;
        RECT  5.770 1.080 6.455 1.240 ;
        RECT  5.730 0.710 5.770 1.700 ;
        RECT  5.650 0.710 5.730 2.080 ;
        RECT  5.170 0.710 5.650 0.870 ;
        RECT  5.570 1.580 5.650 2.080 ;
        RECT  7.715 1.050 7.950 1.270 ;
        RECT  7.595 0.470 7.715 1.270 ;
        RECT  4.660 0.470 7.595 0.590 ;
        RECT  4.660 1.460 5.090 1.620 ;
        RECT  4.500 0.470 4.660 1.620 ;
        RECT  4.020 0.710 4.500 0.870 ;
        RECT  5.010 0.710 5.170 1.290 ;
        RECT  3.690 0.710 3.840 1.440 ;
        RECT  0.750 1.640 0.885 2.060 ;
        RECT  2.010 1.930 2.250 2.090 ;
        RECT  2.320 1.250 2.480 1.700 ;
        RECT  1.800 1.650 2.050 1.810 ;
        RECT  4.190 1.480 4.500 1.620 ;
        RECT  0.060 1.640 0.280 2.060 ;
        LAYER M1 ;
        RECT  6.340 0.760 6.455 0.920 ;
        RECT  6.360 1.650 6.455 2.030 ;
        RECT  7.305 0.760 7.410 0.920 ;
        RECT  7.305 1.650 7.390 2.030 ;
        RECT  7.890 0.490 8.055 0.870 ;
        RECT  7.890 1.650 8.055 2.030 ;
    END
END DFSND4

MACRO DFXD1
    CLASS CORE ;
    FOREIGN DFXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.080 1.940 7.110 2.100 ;
        RECT  7.110 1.390 7.150 2.100 ;
        RECT  7.110 0.420 7.150 0.960 ;
        RECT  7.150 0.420 7.270 2.100 ;
        RECT  7.270 1.940 7.300 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.420 1.540 6.490 2.040 ;
        RECT  6.390 0.710 6.490 0.870 ;
        RECT  6.490 0.710 6.580 2.040 ;
        RECT  6.580 0.710 6.630 1.660 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.960 1.530 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.080 0.790 1.240 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.590 ;
        RECT  0.690 -0.300 1.830 0.300 ;
        RECT  1.830 -0.300 2.050 0.340 ;
        RECT  2.050 -0.300 2.360 0.300 ;
        RECT  2.360 -0.300 2.580 0.340 ;
        RECT  2.580 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.770 ;
        RECT  4.330 -0.300 5.640 0.300 ;
        RECT  5.640 -0.300 5.860 0.340 ;
        RECT  5.860 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.920 0.690 2.820 ;
        RECT  0.690 2.220 1.770 2.820 ;
        RECT  1.770 2.180 1.990 2.820 ;
        RECT  1.990 2.220 2.360 2.820 ;
        RECT  2.360 2.180 2.580 2.820 ;
        RECT  2.580 2.220 4.020 2.820 ;
        RECT  4.020 2.040 4.240 2.820 ;
        RECT  4.240 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.300 1.080 6.370 1.240 ;
        RECT  4.900 0.750 4.990 2.050 ;
        RECT  4.990 0.750 5.040 0.990 ;
        RECT  4.990 1.930 5.780 2.050 ;
        RECT  5.780 1.660 5.900 2.050 ;
        RECT  5.900 1.660 5.920 1.780 ;
        RECT  5.920 1.440 6.060 1.780 ;
        RECT  5.110 1.270 5.160 1.770 ;
        RECT  4.960 0.470 5.160 0.590 ;
        RECT  5.160 0.470 5.240 1.770 ;
        RECT  5.240 0.470 5.280 1.390 ;
        RECT  3.980 1.130 4.100 1.600 ;
        RECT  4.100 1.480 4.450 1.600 ;
        RECT  4.450 1.480 4.560 1.980 ;
        RECT  4.520 0.700 4.560 0.920 ;
        RECT  4.560 0.700 4.610 1.980 ;
        RECT  4.610 0.700 4.680 1.600 ;
        RECT  3.460 0.610 3.580 0.770 ;
        RECT  3.580 0.610 3.700 1.770 ;
        RECT  3.700 0.890 4.280 1.010 ;
        RECT  4.280 0.890 4.400 1.340 ;
        RECT  4.400 1.100 4.440 1.340 ;
        RECT  2.790 0.710 2.950 0.970 ;
        RECT  2.950 0.850 3.070 1.720 ;
        RECT  3.070 1.240 3.460 1.400 ;
        RECT  1.400 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.290 0.730 ;
        RECT  1.310 1.930 3.040 2.050 ;
        RECT  3.040 1.930 3.280 2.090 ;
        RECT  2.050 0.710 2.330 0.870 ;
        RECT  2.330 0.710 2.450 1.810 ;
        RECT  2.450 1.120 2.830 1.290 ;
        RECT  0.070 0.710 0.910 0.870 ;
        RECT  0.910 0.710 1.030 1.800 ;
        RECT  1.030 1.080 1.210 1.240 ;
        RECT  1.030 0.710 1.690 0.830 ;
        RECT  1.690 0.710 1.850 1.030 ;
        RECT  6.260 1.080 6.300 2.060 ;
        RECT  6.180 0.710 6.260 2.060 ;
        RECT  6.140 0.710 6.180 1.240 ;
        RECT  6.020 1.900 6.180 2.060 ;
        RECT  5.780 0.710 6.140 0.860 ;
        RECT  6.990 1.050 7.030 1.290 ;
        RECT  6.870 0.470 6.990 1.290 ;
        RECT  5.520 0.470 6.870 0.590 ;
        RECT  5.400 0.470 5.520 1.810 ;
        RECT  5.360 1.590 5.400 1.810 ;
        RECT  5.640 0.710 5.780 1.400 ;
        RECT  4.850 0.870 4.900 2.050 ;
        RECT  4.740 0.430 4.960 0.590 ;
        RECT  3.860 1.130 3.980 1.290 ;
        RECT  3.420 1.610 3.580 1.770 ;
        RECT  2.740 1.560 2.950 1.720 ;
        RECT  1.160 0.430 1.400 0.590 ;
        RECT  1.150 1.620 1.310 2.050 ;
        RECT  2.050 1.650 2.330 1.810 ;
        RECT  0.070 1.640 0.910 1.800 ;
    END
END DFXD1

MACRO DFXD2
    CLASS CORE ;
    FOREIGN DFXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.310 1.940 8.340 2.100 ;
        RECT  8.340 1.390 8.410 2.100 ;
        RECT  8.340 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.500 2.100 ;
        RECT  8.500 1.940 8.530 2.100 ;
        RECT  8.500 0.780 8.550 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.605 1.940 7.635 2.100 ;
        RECT  7.635 1.390 7.770 2.100 ;
        RECT  7.585 0.710 7.770 0.870 ;
        RECT  7.770 0.710 7.795 2.100 ;
        RECT  7.795 1.940 7.825 2.100 ;
        RECT  7.795 0.710 7.910 1.515 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.835 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 2.040 0.300 ;
        RECT  2.040 -0.300 2.260 0.340 ;
        RECT  2.260 -0.300 2.805 0.300 ;
        RECT  2.805 -0.300 3.025 0.340 ;
        RECT  3.025 -0.300 4.665 0.300 ;
        RECT  4.665 -0.300 4.885 0.340 ;
        RECT  4.885 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.930 2.820 ;
        RECT  1.930 2.180 2.155 2.820 ;
        RECT  2.155 2.220 2.810 2.820 ;
        RECT  2.810 2.180 3.030 2.820 ;
        RECT  3.030 2.220 4.665 2.820 ;
        RECT  4.665 2.020 4.885 2.820 ;
        RECT  4.885 2.220 6.415 2.820 ;
        RECT  6.415 2.180 6.635 2.820 ;
        RECT  6.635 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.395 1.240 3.855 1.400 ;
        RECT  1.440 0.470 3.565 0.590 ;
        RECT  3.565 0.460 3.805 0.620 ;
        RECT  1.340 1.890 3.595 2.010 ;
        RECT  3.595 1.660 3.755 2.010 ;
        RECT  2.490 0.710 3.015 0.870 ;
        RECT  3.015 0.710 3.135 1.770 ;
        RECT  3.135 1.050 3.155 1.270 ;
        RECT  1.600 1.605 1.770 1.770 ;
        RECT  1.600 0.710 1.860 0.870 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 1.030 0.880 ;
        RECT  1.030 0.760 1.190 1.290 ;
        RECT  3.275 0.710 3.395 1.755 ;
        RECT  3.255 0.710 3.275 0.930 ;
        RECT  4.895 1.050 5.055 1.630 ;
        RECT  4.135 1.510 4.895 1.630 ;
        RECT  5.185 0.760 5.310 1.910 ;
        RECT  4.735 0.760 5.185 0.920 ;
        RECT  5.045 1.750 5.185 1.910 ;
        RECT  5.980 1.320 6.025 1.540 ;
        RECT  5.860 0.470 5.980 1.540 ;
        RECT  4.425 0.470 5.860 0.610 ;
        RECT  6.825 1.030 6.985 1.510 ;
        RECT  6.605 1.390 6.825 1.510 ;
        RECT  6.485 1.390 6.605 2.050 ;
        RECT  5.635 1.930 6.485 2.050 ;
        RECT  7.270 1.080 7.650 1.240 ;
        RECT  7.265 0.710 7.270 1.240 ;
        RECT  7.105 0.710 7.265 1.750 ;
        RECT  6.575 0.710 7.105 0.870 ;
        RECT  7.100 1.630 7.105 1.750 ;
        RECT  6.880 1.630 7.100 2.050 ;
        RECT  8.200 1.050 8.270 1.270 ;
        RECT  8.080 0.470 8.200 1.270 ;
        RECT  6.315 0.470 8.080 0.590 ;
        RECT  6.155 0.470 6.315 1.810 ;
        RECT  6.435 0.710 6.575 1.270 ;
        RECT  5.995 1.660 6.155 1.810 ;
        RECT  5.475 0.730 5.635 2.050 ;
        RECT  4.255 0.470 4.425 0.710 ;
        RECT  4.575 0.760 4.735 1.320 ;
        RECT  3.975 0.440 4.135 1.910 ;
        RECT  3.255 1.535 3.275 1.755 ;
        RECT  1.200 0.430 1.440 0.590 ;
        RECT  1.180 1.580 1.340 2.010 ;
        RECT  2.395 1.610 3.015 1.770 ;
        RECT  1.460 0.710 1.600 1.770 ;
        RECT  0.080 0.590 0.200 1.850 ;
    END
END DFXD2

MACRO DFXD4
    CLASS CORE ;
    FOREIGN DFXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.550 1.650 9.870 2.030 ;
        RECT  9.550 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 2.030 ;
        RECT  10.290 1.650 10.460 2.030 ;
        RECT  10.290 0.490 10.460 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.170 1.650 8.590 2.030 ;
        RECT  8.150 0.760 8.590 0.920 ;
        RECT  8.590 0.760 9.010 2.030 ;
        RECT  9.010 1.650 9.080 2.030 ;
        RECT  9.010 0.760 9.100 0.920 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.080 2.010 1.240 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.070 2.745 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 4.560 0.300 ;
        RECT  4.560 -0.300 4.780 0.340 ;
        RECT  4.780 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.930 2.820 ;
        RECT  1.930 2.180 2.155 2.820 ;
        RECT  2.155 2.220 2.710 2.820 ;
        RECT  2.710 2.180 2.930 2.820 ;
        RECT  2.930 2.220 4.560 2.820 ;
        RECT  4.560 2.040 4.780 2.820 ;
        RECT  4.780 2.220 7.080 2.820 ;
        RECT  7.080 2.180 7.300 2.820 ;
        RECT  7.300 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 1.050 0.880 ;
        RECT  1.050 0.760 1.190 1.290 ;
        RECT  1.600 0.710 1.860 0.870 ;
        RECT  1.600 1.605 1.770 1.770 ;
        RECT  2.995 1.050 3.015 1.270 ;
        RECT  2.875 0.710 2.995 1.795 ;
        RECT  2.335 0.710 2.875 0.870 ;
        RECT  3.500 1.640 3.660 2.035 ;
        RECT  1.340 1.915 3.500 2.035 ;
        RECT  3.425 0.460 3.665 0.620 ;
        RECT  1.440 0.470 3.425 0.590 ;
        RECT  3.300 1.240 3.760 1.400 ;
        RECT  3.255 1.240 3.300 1.775 ;
        RECT  3.135 0.710 3.255 1.775 ;
        RECT  4.790 1.050 4.950 1.630 ;
        RECT  4.040 1.510 4.790 1.630 ;
        RECT  3.980 0.990 4.040 1.910 ;
        RECT  3.880 0.460 3.980 1.910 ;
        RECT  5.070 0.770 5.190 1.910 ;
        RECT  4.630 0.770 5.070 0.920 ;
        RECT  4.940 1.750 5.070 1.910 ;
        RECT  5.890 1.320 5.940 1.540 ;
        RECT  5.750 0.470 5.890 1.540 ;
        RECT  4.320 0.470 5.750 0.590 ;
        RECT  7.510 1.030 7.670 1.480 ;
        RECT  7.325 1.360 7.510 1.480 ;
        RECT  7.205 1.360 7.325 2.010 ;
        RECT  5.530 1.890 7.205 2.010 ;
        RECT  7.940 1.080 8.280 1.240 ;
        RECT  7.820 0.710 7.940 1.750 ;
        RECT  7.285 0.710 7.820 0.870 ;
        RECT  7.670 1.600 7.820 1.750 ;
        RECT  7.510 1.600 7.670 2.100 ;
        RECT  7.165 0.710 7.285 1.170 ;
        RECT  6.580 1.050 7.165 1.170 ;
        RECT  9.430 1.080 9.640 1.240 ;
        RECT  9.310 0.470 9.430 1.240 ;
        RECT  6.955 0.470 9.310 0.590 ;
        RECT  6.250 1.610 7.005 1.770 ;
        RECT  6.795 0.470 6.955 0.840 ;
        RECT  6.250 0.650 6.795 0.840 ;
        RECT  6.110 0.650 6.250 1.770 ;
        RECT  6.030 0.650 6.110 0.840 ;
        RECT  6.420 1.050 6.580 1.290 ;
        RECT  6.060 1.540 6.110 1.770 ;
        RECT  5.370 0.710 5.530 2.010 ;
        RECT  4.100 0.430 4.320 0.590 ;
        RECT  4.470 0.770 4.630 1.320 ;
        RECT  3.835 0.460 3.880 1.120 ;
        RECT  3.115 0.710 3.135 0.930 ;
        RECT  1.200 0.430 1.440 0.590 ;
        RECT  1.180 1.580 1.340 2.035 ;
        RECT  2.285 1.635 2.875 1.795 ;
        RECT  1.460 0.710 1.600 1.770 ;
        RECT  0.080 0.590 0.200 1.850 ;
        LAYER M1 ;
        RECT  8.150 0.760 8.375 0.920 ;
        RECT  9.550 0.490 9.655 0.870 ;
        RECT  8.170 1.650 8.375 2.030 ;
        RECT  9.550 1.650 9.655 2.030 ;
    END
END DFXD4

MACRO EDFCND1
    CLASS CORE ;
    FOREIGN EDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.680 1.940 8.710 2.100 ;
        RECT  8.710 1.390 8.730 2.100 ;
        RECT  8.710 0.420 8.730 0.900 ;
        RECT  8.730 0.420 8.870 2.100 ;
        RECT  8.870 1.940 8.900 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.960 1.450 8.090 1.610 ;
        RECT  7.960 0.710 8.090 0.870 ;
        RECT  8.090 0.710 8.230 1.610 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.090 1.005 7.590 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.640 ;
        RECT  7.110 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.600 2.820 ;
        RECT  2.600 2.180 2.820 2.820 ;
        RECT  2.820 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 6.670 2.820 ;
        RECT  6.670 2.180 6.890 2.820 ;
        RECT  6.890 2.220 7.490 2.820 ;
        RECT  7.490 2.180 7.710 2.820 ;
        RECT  7.710 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.010 1.690 3.440 1.810 ;
        RECT  3.440 1.690 3.560 2.050 ;
        RECT  3.560 1.930 4.810 2.050 ;
        RECT  4.810 1.820 4.930 2.050 ;
        RECT  4.930 1.820 5.610 1.940 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.480 0.760 6.520 0.880 ;
        RECT  6.480 1.430 6.600 1.570 ;
        RECT  6.520 0.630 6.680 0.880 ;
        RECT  6.680 0.760 7.265 0.880 ;
        RECT  7.265 0.470 7.385 0.880 ;
        RECT  5.730 1.930 8.370 2.050 ;
        RECT  7.385 0.470 8.370 0.590 ;
        RECT  8.370 0.470 8.510 2.050 ;
        RECT  8.510 1.050 8.610 1.270 ;
        RECT  6.735 1.080 6.855 1.570 ;
        RECT  6.855 1.430 7.720 1.570 ;
        RECT  7.520 0.710 7.720 0.870 ;
        RECT  7.720 0.710 7.840 1.570 ;
        RECT  7.840 1.050 7.970 1.270 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  6.190 1.690 7.870 1.810 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.840 1.800 ;
        RECT  3.840 0.720 3.940 1.200 ;
        RECT  3.940 1.060 4.870 1.200 ;
        RECT  4.870 1.040 5.110 1.200 ;
        RECT  4.570 1.580 4.690 1.810 ;
        RECT  4.690 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.570 ;
        RECT  3.240 1.140 3.560 1.300 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.100 2.050 ;
        RECT  3.100 1.930 3.320 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  6.600 1.080 6.735 1.240 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.680 1.060 3.780 1.800 ;
        RECT  4.020 1.650 4.570 1.810 ;
        RECT  3.000 1.410 3.120 1.570 ;
        RECT  1.290 0.470 1.450 0.740 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
        RECT  1.850 1.360 2.010 1.810 ;
    END
END EDFCND1

MACRO EDFCND2
    CLASS CORE ;
    FOREIGN EDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.270 1.940 9.300 2.100 ;
        RECT  9.300 1.390 9.460 2.100 ;
        RECT  9.300 0.420 9.460 0.900 ;
        RECT  9.460 1.940 9.490 2.100 ;
        RECT  9.460 1.390 9.690 1.515 ;
        RECT  9.460 0.780 9.690 0.900 ;
        RECT  9.690 0.780 9.830 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.590 1.590 8.730 1.810 ;
        RECT  8.590 0.710 8.730 0.930 ;
        RECT  8.730 0.710 8.870 1.810 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 1.285 8.230 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.490 ;
        RECT  7.110 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 1.960 2.820 ;
        RECT  1.960 2.180 2.180 2.820 ;
        RECT  2.180 2.220 2.600 2.820 ;
        RECT  2.600 2.180 2.820 2.820 ;
        RECT  2.820 2.220 4.620 2.820 ;
        RECT  4.620 2.060 4.840 2.820 ;
        RECT  4.840 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.730 1.930 9.030 2.050 ;
        RECT  7.390 0.470 9.030 0.590 ;
        RECT  9.030 0.470 9.150 2.050 ;
        RECT  9.150 1.050 9.250 1.270 ;
        RECT  6.800 0.890 6.920 1.570 ;
        RECT  6.920 1.430 7.290 1.570 ;
        RECT  6.920 0.890 7.540 1.010 ;
        RECT  7.540 0.710 7.760 1.010 ;
        RECT  7.760 1.650 8.350 1.810 ;
        RECT  7.760 0.890 8.350 1.010 ;
        RECT  8.350 0.890 8.470 1.810 ;
        RECT  8.470 1.050 8.600 1.270 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  6.190 1.690 7.410 1.810 ;
        RECT  7.400 1.130 7.410 1.320 ;
        RECT  7.410 1.130 7.530 1.810 ;
        RECT  7.530 1.130 7.620 1.320 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.920 1.570 ;
        RECT  3.920 0.720 3.940 1.200 ;
        RECT  3.940 1.060 4.870 1.200 ;
        RECT  4.870 1.040 5.110 1.200 ;
        RECT  4.260 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.510 ;
        RECT  3.240 1.150 3.580 1.270 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.260 2.050 ;
        RECT  3.260 1.930 3.500 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  7.270 0.470 7.390 0.770 ;
        RECT  6.680 0.650 7.270 0.770 ;
        RECT  6.520 0.650 6.680 0.880 ;
        RECT  6.480 1.430 6.620 1.570 ;
        RECT  6.480 0.760 6.520 0.880 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  4.500 1.820 5.610 1.940 ;
        RECT  4.380 1.820 4.500 2.050 ;
        RECT  3.920 1.930 4.380 2.050 ;
        RECT  3.800 1.690 3.920 2.050 ;
        RECT  1.980 1.690 3.800 1.810 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  6.600 1.080 6.800 1.240 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.630 1.410 3.780 1.570 ;
        RECT  4.040 1.580 4.260 1.740 ;
        RECT  3.000 1.350 3.120 1.510 ;
        RECT  1.290 0.470 1.450 0.710 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFCND2

MACRO EDFCND4
    CLASS CORE ;
    FOREIGN EDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.510 1.650 10.830 2.030 ;
        RECT  10.510 0.490 10.830 0.870 ;
        RECT  10.830 0.490 11.250 2.030 ;
        RECT  11.250 1.650 11.420 2.030 ;
        RECT  11.250 0.490 11.420 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.110 1.600 9.230 1.760 ;
        RECT  9.110 0.760 9.230 0.920 ;
        RECT  9.230 0.760 9.650 1.760 ;
        RECT  9.650 1.600 10.060 1.760 ;
        RECT  9.650 0.760 10.060 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.090 1.005 8.550 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.490 ;
        RECT  7.110 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 4.620 2.820 ;
        RECT  4.620 2.060 4.840 2.820 ;
        RECT  4.840 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.920 1.570 ;
        RECT  3.920 0.720 3.940 1.200 ;
        RECT  3.940 1.060 4.870 1.200 ;
        RECT  4.870 1.040 5.110 1.200 ;
        RECT  4.040 1.580 4.260 1.740 ;
        RECT  4.260 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.510 ;
        RECT  3.240 1.150 3.580 1.270 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.260 2.050 ;
        RECT  3.260 1.930 3.500 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  7.420 1.100 7.580 1.810 ;
        RECT  6.190 1.690 7.420 1.810 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  8.700 1.030 8.860 1.630 ;
        RECT  7.900 1.470 8.700 1.630 ;
        RECT  7.780 0.850 7.900 1.630 ;
        RECT  7.730 0.850 7.780 0.970 ;
        RECT  7.570 0.720 7.730 0.970 ;
        RECT  7.075 0.850 7.570 0.970 ;
        RECT  7.075 1.430 7.290 1.570 ;
        RECT  6.955 0.850 7.075 1.570 ;
        RECT  10.360 1.080 10.615 1.240 ;
        RECT  10.240 0.470 10.360 2.050 ;
        RECT  7.390 0.470 10.240 0.590 ;
        RECT  5.730 1.930 10.240 2.050 ;
        RECT  7.270 0.470 7.390 0.730 ;
        RECT  6.680 0.610 7.270 0.730 ;
        RECT  6.520 0.610 6.680 0.880 ;
        RECT  6.480 1.430 6.620 1.570 ;
        RECT  6.480 0.760 6.520 0.880 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  4.500 1.820 5.610 1.940 ;
        RECT  4.380 1.820 4.500 2.050 ;
        RECT  3.920 1.930 4.380 2.050 ;
        RECT  3.800 1.690 3.920 2.050 ;
        RECT  1.980 1.690 3.800 1.810 ;
        RECT  6.600 1.080 6.955 1.240 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.630 1.410 3.780 1.570 ;
        RECT  3.000 1.350 3.120 1.510 ;
        RECT  1.290 0.470 1.450 0.710 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
        LAYER M1 ;
        RECT  10.510 1.650 10.615 2.030 ;
        RECT  10.510 0.490 10.615 0.870 ;
        RECT  9.865 1.600 10.060 1.760 ;
        RECT  9.865 0.760 10.060 0.920 ;
    END
END EDFCND4

MACRO EDFCNQD1
    CLASS CORE ;
    FOREIGN EDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.960 1.450 8.090 1.610 ;
        RECT  7.960 0.710 8.090 0.870 ;
        RECT  8.090 0.710 8.230 1.610 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.090 1.005 7.590 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.910 0.300 ;
        RECT  1.910 -0.300 2.130 0.340 ;
        RECT  2.130 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.640 ;
        RECT  7.110 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.600 2.820 ;
        RECT  2.600 2.180 2.820 2.820 ;
        RECT  2.820 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 6.670 2.820 ;
        RECT  6.670 2.180 6.890 2.820 ;
        RECT  6.890 2.220 7.490 2.820 ;
        RECT  7.490 2.180 7.710 2.820 ;
        RECT  7.710 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.930 1.820 5.610 1.940 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.480 0.760 6.520 0.880 ;
        RECT  6.480 1.430 6.600 1.570 ;
        RECT  6.520 0.630 6.680 0.880 ;
        RECT  6.680 0.760 7.265 0.880 ;
        RECT  7.265 0.470 7.385 0.880 ;
        RECT  5.730 1.930 8.350 2.050 ;
        RECT  7.385 0.470 8.350 0.590 ;
        RECT  8.350 0.470 8.470 2.050 ;
        RECT  6.735 1.080 6.855 1.570 ;
        RECT  6.855 1.430 7.720 1.570 ;
        RECT  7.520 0.710 7.720 0.870 ;
        RECT  7.720 0.710 7.840 1.570 ;
        RECT  7.840 1.050 7.970 1.270 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  6.190 1.690 7.870 1.810 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.840 1.800 ;
        RECT  3.840 0.720 3.940 1.200 ;
        RECT  3.940 1.060 4.870 1.200 ;
        RECT  4.870 1.040 5.110 1.200 ;
        RECT  4.570 1.580 4.690 1.810 ;
        RECT  4.690 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.570 ;
        RECT  3.240 1.140 3.560 1.300 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.100 2.050 ;
        RECT  3.100 1.930 3.320 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  4.810 1.820 4.930 2.050 ;
        RECT  3.560 1.930 4.810 2.050 ;
        RECT  3.440 1.690 3.560 2.050 ;
        RECT  2.010 1.690 3.440 1.810 ;
        RECT  1.850 1.360 2.010 1.810 ;
        RECT  6.600 1.080 6.735 1.240 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.680 1.060 3.780 1.800 ;
        RECT  4.020 1.650 4.570 1.810 ;
        RECT  3.000 1.410 3.120 1.570 ;
        RECT  1.290 0.470 1.450 0.740 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFCNQD1

MACRO EDFCNQD2
    CLASS CORE ;
    FOREIGN EDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.590 1.590 8.730 1.810 ;
        RECT  8.590 0.710 8.730 0.930 ;
        RECT  8.730 0.710 8.870 1.810 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 1.285 8.230 1.520 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.490 ;
        RECT  7.110 -0.300 8.940 0.300 ;
        RECT  8.940 -0.300 9.160 0.340 ;
        RECT  9.160 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 1.960 2.820 ;
        RECT  1.960 2.180 2.180 2.820 ;
        RECT  2.180 2.220 2.600 2.820 ;
        RECT  2.600 2.180 2.820 2.820 ;
        RECT  2.820 2.220 4.620 2.820 ;
        RECT  4.620 2.060 4.840 2.820 ;
        RECT  4.840 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 6.670 2.820 ;
        RECT  6.670 2.180 6.890 2.820 ;
        RECT  6.890 2.220 8.940 2.820 ;
        RECT  8.940 2.180 9.160 2.820 ;
        RECT  9.160 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.680 0.650 7.270 0.770 ;
        RECT  7.270 0.470 7.390 0.770 ;
        RECT  5.730 1.930 9.030 2.050 ;
        RECT  7.390 0.470 9.030 0.590 ;
        RECT  9.030 0.470 9.150 2.050 ;
        RECT  6.800 0.890 6.920 1.570 ;
        RECT  6.920 1.430 7.310 1.570 ;
        RECT  6.920 0.890 7.540 1.010 ;
        RECT  7.540 0.750 7.760 1.010 ;
        RECT  7.760 1.650 8.350 1.810 ;
        RECT  7.760 0.890 8.350 1.010 ;
        RECT  8.350 0.890 8.470 1.810 ;
        RECT  8.470 1.050 8.600 1.270 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  6.190 1.690 7.500 1.810 ;
        RECT  7.380 1.150 7.500 1.310 ;
        RECT  7.500 1.150 7.620 1.810 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.920 1.570 ;
        RECT  3.920 0.720 3.940 1.180 ;
        RECT  3.940 1.040 5.110 1.180 ;
        RECT  4.260 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.510 ;
        RECT  3.240 1.130 3.580 1.290 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.260 2.050 ;
        RECT  3.260 1.930 3.500 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  6.530 0.650 6.680 0.880 ;
        RECT  6.480 1.430 6.620 1.570 ;
        RECT  6.480 0.760 6.530 0.880 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  4.500 1.820 5.610 1.940 ;
        RECT  4.380 1.820 4.500 2.050 ;
        RECT  3.920 1.930 4.380 2.050 ;
        RECT  3.800 1.690 3.920 2.050 ;
        RECT  1.990 1.690 3.800 1.810 ;
        RECT  6.600 1.080 6.800 1.240 ;
        RECT  1.830 1.360 1.990 1.810 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.630 1.410 3.780 1.570 ;
        RECT  4.040 1.580 4.260 1.740 ;
        RECT  3.000 1.350 3.120 1.510 ;
        RECT  1.290 0.470 1.450 0.710 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFCNQD2

MACRO EDFCNQD4
    CLASS CORE ;
    FOREIGN EDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.590 1.650 8.910 1.810 ;
        RECT  8.570 0.760 8.910 0.920 ;
        RECT  8.910 0.760 9.330 1.810 ;
        RECT  9.330 1.650 9.500 1.810 ;
        RECT  9.330 0.760 9.500 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.050 0.990 8.090 1.230 ;
        RECT  8.090 0.990 8.230 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 4.650 0.300 ;
        RECT  4.650 -0.300 4.880 0.680 ;
        RECT  4.880 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.490 ;
        RECT  7.110 -0.300 8.180 0.300 ;
        RECT  8.180 -0.300 8.400 0.340 ;
        RECT  8.400 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 4.620 2.820 ;
        RECT  4.620 2.060 4.840 2.820 ;
        RECT  4.840 2.220 5.220 2.820 ;
        RECT  5.220 2.060 5.440 2.820 ;
        RECT  5.440 2.220 6.670 2.820 ;
        RECT  6.670 2.180 6.890 2.820 ;
        RECT  6.890 2.220 8.180 2.820 ;
        RECT  8.180 2.180 8.400 2.820 ;
        RECT  8.400 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.955 0.890 7.075 1.570 ;
        RECT  7.075 1.430 7.310 1.570 ;
        RECT  7.075 0.890 7.540 1.010 ;
        RECT  7.540 0.710 7.760 1.010 ;
        RECT  7.780 1.650 7.810 1.810 ;
        RECT  7.760 0.890 7.810 1.010 ;
        RECT  7.810 0.890 7.930 1.810 ;
        RECT  7.930 1.650 8.350 1.810 ;
        RECT  8.350 1.080 8.470 1.810 ;
        RECT  8.470 1.080 8.695 1.240 ;
        RECT  5.760 1.300 6.030 1.420 ;
        RECT  6.030 1.300 6.190 1.810 ;
        RECT  6.190 1.690 7.490 1.810 ;
        RECT  7.370 1.150 7.490 1.310 ;
        RECT  7.490 1.150 7.610 1.810 ;
        RECT  4.130 0.440 4.250 0.920 ;
        RECT  4.250 0.800 5.000 0.920 ;
        RECT  5.000 0.470 5.120 0.920 ;
        RECT  5.120 0.470 6.180 0.590 ;
        RECT  6.180 0.470 6.400 0.630 ;
        RECT  5.240 0.710 5.380 1.700 ;
        RECT  5.380 1.540 5.860 1.700 ;
        RECT  3.780 0.720 3.920 1.570 ;
        RECT  3.920 0.720 3.940 1.200 ;
        RECT  3.940 1.060 4.870 1.200 ;
        RECT  4.870 1.040 5.110 1.200 ;
        RECT  4.260 1.580 4.950 1.700 ;
        RECT  3.000 0.710 3.120 0.850 ;
        RECT  3.120 0.710 3.240 1.510 ;
        RECT  3.240 1.150 3.580 1.270 ;
        RECT  1.450 0.470 3.380 0.590 ;
        RECT  3.380 0.470 3.540 0.730 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.260 2.050 ;
        RECT  3.260 1.930 3.500 2.090 ;
        RECT  2.280 0.710 2.760 0.850 ;
        RECT  2.760 0.710 2.880 1.510 ;
        RECT  2.880 1.020 2.990 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  9.620 0.470 9.740 2.050 ;
        RECT  7.390 0.470 9.620 0.590 ;
        RECT  5.730 1.930 9.620 2.050 ;
        RECT  7.270 0.470 7.390 0.770 ;
        RECT  6.690 0.650 7.270 0.770 ;
        RECT  6.530 0.650 6.690 0.880 ;
        RECT  6.480 1.430 6.620 1.570 ;
        RECT  6.480 0.760 6.530 0.880 ;
        RECT  6.360 0.760 6.480 1.570 ;
        RECT  6.060 0.760 6.360 0.920 ;
        RECT  5.610 1.820 5.730 2.050 ;
        RECT  4.500 1.820 5.610 1.940 ;
        RECT  4.380 1.820 4.500 2.050 ;
        RECT  3.920 1.930 4.380 2.050 ;
        RECT  3.800 1.690 3.920 2.050 ;
        RECT  1.980 1.690 3.800 1.810 ;
        RECT  6.600 1.080 6.955 1.240 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  5.600 0.710 5.760 1.420 ;
        RECT  3.920 0.440 4.130 0.600 ;
        RECT  4.220 1.320 5.240 1.460 ;
        RECT  3.630 1.410 3.780 1.570 ;
        RECT  4.040 1.580 4.260 1.740 ;
        RECT  3.000 1.350 3.120 1.510 ;
        RECT  1.290 0.470 1.450 0.710 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  2.280 1.355 2.760 1.510 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
        LAYER M1 ;
        RECT  8.590 1.650 8.695 1.810 ;
        RECT  8.570 0.760 8.695 0.920 ;
    END
END EDFCNQD4

MACRO EDFD1
    CLASS CORE ;
    FOREIGN EDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.400 1.960 7.430 2.100 ;
        RECT  7.430 0.420 7.590 2.100 ;
        RECT  7.590 1.960 7.620 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.600 1.410 6.810 1.810 ;
        RECT  6.600 0.710 6.810 0.870 ;
        RECT  6.810 0.710 6.820 1.810 ;
        RECT  6.820 0.710 6.950 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.910 0.300 ;
        RECT  1.910 -0.300 2.130 0.340 ;
        RECT  2.130 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.720 ;
        RECT  4.580 -0.300 7.000 0.300 ;
        RECT  7.000 -0.300 7.220 0.340 ;
        RECT  7.220 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.280 2.820 ;
        RECT  4.280 1.970 4.500 2.820 ;
        RECT  4.500 2.220 7.000 2.820 ;
        RECT  7.000 2.180 7.220 2.820 ;
        RECT  7.220 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.940 1.020 6.350 1.140 ;
        RECT  6.230 0.710 6.350 0.850 ;
        RECT  6.350 0.710 6.470 1.810 ;
        RECT  6.470 1.080 6.690 1.240 ;
        RECT  5.320 0.470 5.440 1.070 ;
        RECT  5.030 1.690 5.540 1.810 ;
        RECT  5.440 0.950 5.540 1.070 ;
        RECT  5.540 0.950 5.660 1.810 ;
        RECT  5.660 1.310 6.210 1.470 ;
        RECT  5.200 1.270 5.260 1.390 ;
        RECT  5.260 1.270 5.420 1.570 ;
        RECT  4.310 1.420 4.810 1.560 ;
        RECT  4.810 0.445 4.940 1.560 ;
        RECT  3.810 0.840 4.550 0.960 ;
        RECT  4.550 0.840 4.690 1.260 ;
        RECT  2.910 1.410 3.020 1.570 ;
        RECT  2.890 0.710 3.020 0.850 ;
        RECT  3.020 0.710 3.140 1.570 ;
        RECT  3.140 1.080 3.150 1.570 ;
        RECT  3.150 1.080 3.530 1.240 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.230 2.050 ;
        RECT  3.230 1.930 3.470 2.090 ;
        RECT  3.260 0.470 3.420 0.710 ;
        RECT  2.170 0.710 2.650 0.850 ;
        RECT  2.650 0.710 2.770 1.500 ;
        RECT  2.770 1.020 2.900 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  6.230 1.650 6.350 1.810 ;
        RECT  7.120 0.470 7.280 2.050 ;
        RECT  5.740 0.470 7.120 0.590 ;
        RECT  5.690 1.930 7.120 2.050 ;
        RECT  5.580 0.470 5.740 0.740 ;
        RECT  5.470 1.930 5.690 2.090 ;
        RECT  4.850 1.930 5.470 2.050 ;
        RECT  4.730 1.690 4.850 2.050 ;
        RECT  2.050 1.690 4.730 1.810 ;
        RECT  1.900 1.360 2.050 1.810 ;
        RECT  5.780 0.900 5.940 1.140 ;
        RECT  5.160 0.470 5.320 0.630 ;
        RECT  5.060 0.750 5.200 1.390 ;
        RECT  4.150 1.080 4.310 1.560 ;
        RECT  3.650 0.530 3.810 1.570 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.260 0.590 ;
        RECT  2.170 1.360 2.650 1.500 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFD1

MACRO EDFD2
    CLASS CORE ;
    FOREIGN EDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.710 1.390 7.770 1.890 ;
        RECT  7.710 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.870 1.890 ;
        RECT  7.870 0.780 7.910 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.940 1.410 7.130 1.810 ;
        RECT  6.920 0.710 7.130 0.870 ;
        RECT  7.130 0.710 7.160 1.810 ;
        RECT  7.160 0.710 7.270 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.910 0.300 ;
        RECT  1.910 -0.300 2.130 0.340 ;
        RECT  2.130 -0.300 2.480 0.300 ;
        RECT  2.480 -0.300 2.700 0.340 ;
        RECT  2.700 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.720 ;
        RECT  4.580 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 1.960 2.820 ;
        RECT  1.960 2.180 2.180 2.820 ;
        RECT  2.180 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.280 2.820 ;
        RECT  4.280 1.970 4.500 2.820 ;
        RECT  4.500 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.660 1.390 6.250 1.510 ;
        RECT  6.250 1.030 6.410 1.510 ;
        RECT  5.200 1.270 5.260 1.390 ;
        RECT  5.260 1.270 5.420 1.570 ;
        RECT  4.310 1.420 4.810 1.560 ;
        RECT  4.810 0.445 4.940 1.560 ;
        RECT  3.650 0.530 3.810 1.560 ;
        RECT  3.810 1.400 3.840 1.560 ;
        RECT  3.810 0.840 4.550 0.960 ;
        RECT  4.550 0.840 4.690 1.260 ;
        RECT  2.910 1.410 3.020 1.570 ;
        RECT  2.890 0.710 3.020 0.850 ;
        RECT  3.020 0.710 3.140 1.570 ;
        RECT  3.140 1.080 3.150 1.570 ;
        RECT  3.150 1.080 3.530 1.240 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.230 2.050 ;
        RECT  3.230 1.930 3.470 2.090 ;
        RECT  3.260 0.470 3.420 0.710 ;
        RECT  2.170 0.710 2.650 0.850 ;
        RECT  2.650 0.710 2.770 1.560 ;
        RECT  2.770 1.080 2.900 1.240 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  5.540 0.950 5.660 1.810 ;
        RECT  5.440 0.950 5.540 1.070 ;
        RECT  5.030 1.690 5.540 1.810 ;
        RECT  5.320 0.470 5.440 1.070 ;
        RECT  6.745 1.080 6.965 1.240 ;
        RECT  6.625 0.710 6.745 1.810 ;
        RECT  6.040 0.710 6.625 0.850 ;
        RECT  6.230 1.650 6.625 1.810 ;
        RECT  5.940 0.710 6.040 1.170 ;
        RECT  5.920 0.710 5.940 1.270 ;
        RECT  7.440 0.470 7.580 2.050 ;
        RECT  5.740 0.470 7.440 0.590 ;
        RECT  5.690 1.930 7.440 2.050 ;
        RECT  5.580 0.470 5.740 0.740 ;
        RECT  5.470 1.930 5.690 2.090 ;
        RECT  4.850 1.930 5.470 2.050 ;
        RECT  4.730 1.690 4.850 2.050 ;
        RECT  1.980 1.690 4.730 1.810 ;
        RECT  5.780 1.050 5.920 1.270 ;
        RECT  5.160 0.470 5.320 0.630 ;
        RECT  5.060 0.750 5.200 1.390 ;
        RECT  4.150 1.080 4.310 1.560 ;
        RECT  3.620 1.400 3.650 1.560 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.260 0.590 ;
        RECT  2.190 1.420 2.650 1.560 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFD2

MACRO EDFD4
    CLASS CORE ;
    FOREIGN EDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.910 1.650 9.230 2.030 ;
        RECT  8.910 0.490 9.230 0.870 ;
        RECT  9.230 0.490 9.650 2.030 ;
        RECT  9.650 1.650 9.820 2.030 ;
        RECT  9.650 0.490 9.820 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.510 1.605 7.950 1.765 ;
        RECT  7.510 0.710 7.950 0.870 ;
        RECT  7.950 0.710 8.370 1.765 ;
        RECT  8.370 1.605 8.460 1.765 ;
        RECT  8.370 0.710 8.460 0.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 4.280 0.300 ;
        RECT  4.280 -0.300 4.500 0.720 ;
        RECT  4.500 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 4.280 2.820 ;
        RECT  4.280 1.970 4.500 2.820 ;
        RECT  4.500 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  2.770 1.080 2.900 1.240 ;
        RECT  2.650 0.710 2.770 1.560 ;
        RECT  2.170 0.710 2.650 0.850 ;
        RECT  3.260 0.470 3.420 0.710 ;
        RECT  3.230 1.930 3.470 2.090 ;
        RECT  1.500 1.930 3.230 2.050 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  3.150 1.080 3.530 1.240 ;
        RECT  3.140 1.080 3.150 1.570 ;
        RECT  3.020 0.710 3.140 1.570 ;
        RECT  2.890 0.710 3.020 0.850 ;
        RECT  4.470 0.840 4.610 1.260 ;
        RECT  3.810 0.840 4.470 0.960 ;
        RECT  3.810 1.400 3.840 1.560 ;
        RECT  3.650 0.530 3.810 1.560 ;
        RECT  4.870 1.425 4.890 1.560 ;
        RECT  4.730 0.540 4.870 1.560 ;
        RECT  4.310 1.420 4.730 1.560 ;
        RECT  6.840 1.030 7.000 1.510 ;
        RECT  5.660 1.390 6.840 1.510 ;
        RECT  5.540 0.950 5.660 1.810 ;
        RECT  5.250 0.950 5.540 1.070 ;
        RECT  5.030 1.650 5.540 1.810 ;
        RECT  7.335 1.080 7.555 1.240 ;
        RECT  7.215 0.730 7.335 1.810 ;
        RECT  6.430 0.730 7.215 0.850 ;
        RECT  6.820 1.650 7.215 1.810 ;
        RECT  6.310 0.730 6.430 1.240 ;
        RECT  8.790 1.080 8.930 1.240 ;
        RECT  8.650 0.470 8.790 2.050 ;
        RECT  5.630 0.470 8.650 0.590 ;
        RECT  6.370 1.930 8.650 2.050 ;
        RECT  6.150 1.670 6.370 2.090 ;
        RECT  5.690 1.930 6.150 2.050 ;
        RECT  5.470 1.930 5.690 2.090 ;
        RECT  5.470 0.470 5.630 0.800 ;
        RECT  4.850 1.930 5.470 2.050 ;
        RECT  4.730 1.690 4.850 2.050 ;
        RECT  1.980 1.690 4.730 1.810 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  6.190 1.080 6.310 1.240 ;
        RECT  5.090 0.540 5.250 1.070 ;
        RECT  4.150 1.080 4.310 1.560 ;
        RECT  3.620 1.400 3.650 1.560 ;
        RECT  2.910 1.410 3.020 1.570 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.260 0.590 ;
        RECT  2.190 1.420 2.650 1.560 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
        LAYER M1 ;
        RECT  8.910 1.650 9.015 2.030 ;
        RECT  8.910 0.490 9.015 0.870 ;
        RECT  7.510 1.605 7.735 1.765 ;
        RECT  7.510 0.710 7.735 0.870 ;
    END
END EDFD4

MACRO EDFKCND1
    CLASS CORE ;
    FOREIGN EDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.400 1.960 7.430 2.100 ;
        RECT  7.430 1.390 7.450 2.100 ;
        RECT  7.430 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.590 2.100 ;
        RECT  7.590 1.960 7.620 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.690 1.410 6.810 1.810 ;
        RECT  6.690 0.710 6.810 0.870 ;
        RECT  6.810 0.710 6.910 1.810 ;
        RECT  6.910 0.710 6.950 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 2.230 0.300 ;
        RECT  2.230 -0.300 2.450 0.340 ;
        RECT  2.450 -0.300 2.760 0.300 ;
        RECT  2.760 -0.300 2.980 0.340 ;
        RECT  2.980 -0.300 4.430 0.300 ;
        RECT  4.430 -0.300 4.650 0.480 ;
        RECT  4.650 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 2.760 2.820 ;
        RECT  2.760 2.180 2.980 2.820 ;
        RECT  2.980 2.220 4.430 2.820 ;
        RECT  4.430 1.960 4.650 2.820 ;
        RECT  4.650 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.890 1.690 4.830 1.810 ;
        RECT  4.830 1.690 4.950 2.050 ;
        RECT  4.950 1.930 5.610 2.050 ;
        RECT  5.610 1.930 5.830 2.090 ;
        RECT  5.690 0.470 5.830 0.710 ;
        RECT  5.830 1.930 7.160 2.050 ;
        RECT  5.830 0.470 7.160 0.590 ;
        RECT  7.160 0.470 7.280 2.050 ;
        RECT  7.280 1.050 7.330 1.270 ;
        RECT  6.310 1.650 6.450 1.810 ;
        RECT  6.340 0.710 6.450 0.990 ;
        RECT  6.450 0.710 6.560 1.810 ;
        RECT  6.560 0.830 6.570 1.810 ;
        RECT  6.570 1.080 6.690 1.240 ;
        RECT  5.450 0.450 5.570 1.240 ;
        RECT  5.190 1.650 5.800 1.810 ;
        RECT  5.570 1.120 5.800 1.240 ;
        RECT  5.800 1.120 5.920 1.810 ;
        RECT  5.920 1.120 6.320 1.280 ;
        RECT  5.330 1.360 5.680 1.520 ;
        RECT  4.550 1.410 4.970 1.570 ;
        RECT  4.810 0.580 4.970 0.740 ;
        RECT  4.970 0.580 5.090 1.570 ;
        RECT  3.910 0.530 4.070 1.570 ;
        RECT  4.070 0.860 4.710 0.980 ;
        RECT  4.710 0.860 4.850 1.290 ;
        RECT  1.450 0.470 3.500 0.590 ;
        RECT  3.500 0.430 3.740 0.590 ;
        RECT  3.160 0.710 3.550 0.860 ;
        RECT  3.550 0.710 3.710 1.570 ;
        RECT  1.360 1.930 2.210 2.050 ;
        RECT  2.210 1.930 2.430 2.090 ;
        RECT  2.430 1.930 3.430 2.050 ;
        RECT  3.430 1.930 3.670 2.090 ;
        RECT  2.450 0.710 2.920 0.860 ;
        RECT  2.920 0.710 3.040 1.570 ;
        RECT  3.040 1.030 3.180 1.190 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  5.770 0.830 6.340 0.990 ;
        RECT  5.230 0.450 5.450 0.610 ;
        RECT  5.210 0.730 5.330 1.520 ;
        RECT  4.390 1.100 4.550 1.570 ;
        RECT  3.830 1.410 3.910 1.570 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  3.160 1.410 3.550 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.450 1.410 2.920 1.570 ;
        RECT  0.190 1.510 0.350 1.900 ;
        RECT  1.730 1.230 1.890 1.810 ;
    END
END EDFKCND1

MACRO EDFKCND2
    CLASS CORE ;
    FOREIGN EDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.975 1.940 8.005 2.100 ;
        RECT  8.005 1.390 8.090 2.100 ;
        RECT  8.005 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.165 2.100 ;
        RECT  8.165 1.940 8.195 2.100 ;
        RECT  8.165 0.780 8.230 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.175 1.410 7.395 1.810 ;
        RECT  7.395 1.410 7.450 1.530 ;
        RECT  7.155 0.710 7.450 0.870 ;
        RECT  7.450 0.710 7.590 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.885 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 2.230 0.300 ;
        RECT  2.230 -0.300 2.450 0.340 ;
        RECT  2.450 -0.300 2.855 0.300 ;
        RECT  2.855 -0.300 3.075 0.340 ;
        RECT  3.075 -0.300 4.545 0.300 ;
        RECT  4.545 -0.300 4.765 0.480 ;
        RECT  4.765 -0.300 7.575 0.300 ;
        RECT  7.575 -0.300 7.795 0.340 ;
        RECT  7.795 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 2.855 2.820 ;
        RECT  2.855 2.180 3.075 2.820 ;
        RECT  3.075 2.220 4.545 2.820 ;
        RECT  4.545 2.040 4.765 2.820 ;
        RECT  4.765 2.220 7.575 2.820 ;
        RECT  7.575 2.180 7.795 2.820 ;
        RECT  7.795 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.645 0.710 3.805 1.570 ;
        RECT  1.360 1.930 2.210 2.050 ;
        RECT  2.210 1.930 2.430 2.090 ;
        RECT  2.430 1.930 3.525 2.050 ;
        RECT  3.525 1.930 3.765 2.090 ;
        RECT  2.545 0.710 3.015 0.860 ;
        RECT  3.015 0.710 3.135 1.570 ;
        RECT  3.135 1.030 3.275 1.190 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  3.255 0.710 3.645 0.860 ;
        RECT  3.595 0.430 3.835 0.590 ;
        RECT  1.450 0.470 3.595 0.590 ;
        RECT  4.825 0.860 4.965 1.290 ;
        RECT  4.185 0.860 4.825 0.980 ;
        RECT  4.025 0.530 4.185 1.570 ;
        RECT  5.085 0.580 5.205 1.570 ;
        RECT  4.925 0.580 5.085 0.740 ;
        RECT  4.665 1.410 5.085 1.570 ;
        RECT  5.445 1.410 5.795 1.550 ;
        RECT  6.035 1.140 6.445 1.280 ;
        RECT  5.915 1.140 6.035 1.810 ;
        RECT  5.685 1.140 5.915 1.260 ;
        RECT  5.305 1.680 5.915 1.810 ;
        RECT  5.565 0.450 5.685 1.260 ;
        RECT  6.695 1.080 7.215 1.240 ;
        RECT  6.575 0.710 6.695 1.810 ;
        RECT  6.465 0.710 6.575 1.010 ;
        RECT  6.455 1.400 6.575 1.810 ;
        RECT  7.850 1.080 7.950 1.240 ;
        RECT  7.710 0.470 7.850 2.050 ;
        RECT  5.945 0.470 7.710 0.590 ;
        RECT  5.945 1.930 7.710 2.050 ;
        RECT  5.805 0.470 5.945 0.710 ;
        RECT  5.725 1.930 5.945 2.090 ;
        RECT  5.065 1.930 5.725 2.050 ;
        RECT  4.945 1.690 5.065 2.050 ;
        RECT  1.890 1.690 4.945 1.810 ;
        RECT  5.875 0.885 6.465 1.010 ;
        RECT  5.325 0.450 5.565 0.610 ;
        RECT  5.325 0.740 5.445 1.550 ;
        RECT  4.505 1.100 4.665 1.570 ;
        RECT  3.945 1.410 4.025 1.570 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  3.255 1.410 3.645 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.545 1.410 3.015 1.570 ;
        RECT  0.190 1.510 0.350 1.900 ;
        RECT  1.730 1.230 1.890 1.810 ;
    END
END EDFKCND2

MACRO EDFKCND4
    CLASS CORE ;
    FOREIGN EDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.195 1.650 9.550 2.030 ;
        RECT  9.195 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 2.030 ;
        RECT  9.970 1.650 10.140 2.030 ;
        RECT  9.970 0.490 10.140 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.685 1.580 7.950 1.740 ;
        RECT  7.685 0.760 7.950 0.920 ;
        RECT  7.950 0.760 8.370 1.740 ;
        RECT  8.370 1.580 8.635 1.740 ;
        RECT  8.370 0.760 8.635 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 4.445 0.300 ;
        RECT  4.445 -0.300 4.665 0.480 ;
        RECT  4.665 -0.300 8.795 0.300 ;
        RECT  8.795 -0.300 9.015 0.340 ;
        RECT  9.015 -0.300 10.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 4.445 2.820 ;
        RECT  4.445 2.040 4.665 2.820 ;
        RECT  4.665 2.220 6.595 2.820 ;
        RECT  6.595 2.180 6.815 2.820 ;
        RECT  6.815 2.220 8.795 2.820 ;
        RECT  8.795 2.180 9.015 2.820 ;
        RECT  9.015 2.220 10.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  3.050 1.030 3.190 1.190 ;
        RECT  2.930 0.710 3.050 1.560 ;
        RECT  2.460 0.710 2.930 0.860 ;
        RECT  3.440 1.930 3.680 2.090 ;
        RECT  2.440 1.930 3.440 2.050 ;
        RECT  2.220 1.930 2.440 2.090 ;
        RECT  1.360 1.930 2.220 2.050 ;
        RECT  3.560 0.710 3.720 1.570 ;
        RECT  3.170 0.710 3.560 0.860 ;
        RECT  3.510 0.430 3.750 0.590 ;
        RECT  1.450 0.470 3.510 0.590 ;
        RECT  4.725 0.860 4.865 1.290 ;
        RECT  4.080 0.860 4.725 0.980 ;
        RECT  3.920 0.430 4.080 1.570 ;
        RECT  4.985 0.580 5.105 1.570 ;
        RECT  4.825 0.580 4.985 0.740 ;
        RECT  4.565 1.410 4.985 1.570 ;
        RECT  5.345 1.380 5.695 1.520 ;
        RECT  5.935 1.140 6.985 1.260 ;
        RECT  5.815 1.140 5.935 1.810 ;
        RECT  5.585 1.140 5.815 1.260 ;
        RECT  5.205 1.650 5.815 1.810 ;
        RECT  5.465 0.450 5.585 1.260 ;
        RECT  7.255 1.050 7.735 1.270 ;
        RECT  7.225 0.830 7.255 1.810 ;
        RECT  7.115 0.710 7.225 1.810 ;
        RECT  6.995 0.710 7.115 1.020 ;
        RECT  6.975 1.650 7.115 1.810 ;
        RECT  8.975 1.080 9.305 1.240 ;
        RECT  8.855 0.470 8.975 2.050 ;
        RECT  5.845 0.470 8.855 0.590 ;
        RECT  6.555 1.930 8.855 2.050 ;
        RECT  6.335 1.725 6.555 2.050 ;
        RECT  5.845 1.930 6.335 2.050 ;
        RECT  5.705 0.470 5.845 0.710 ;
        RECT  5.625 1.930 5.845 2.090 ;
        RECT  4.965 1.930 5.625 2.050 ;
        RECT  4.845 1.690 4.965 2.050 ;
        RECT  1.890 1.690 4.845 1.810 ;
        RECT  1.730 1.230 1.890 1.810 ;
        RECT  5.990 0.880 6.995 1.020 ;
        RECT  5.245 0.450 5.465 0.610 ;
        RECT  5.225 0.730 5.345 1.520 ;
        RECT  4.405 1.100 4.565 1.570 ;
        RECT  3.840 1.410 3.920 1.570 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  3.170 1.410 3.560 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.460 1.400 2.930 1.560 ;
        RECT  0.190 1.510 0.350 1.900 ;
        LAYER M1 ;
        RECT  9.195 1.650 9.335 2.030 ;
        RECT  9.195 0.490 9.335 0.870 ;
        RECT  8.585 1.580 8.635 1.740 ;
        RECT  8.585 0.760 8.635 0.920 ;
        RECT  7.685 1.580 7.735 1.740 ;
        RECT  7.685 0.760 7.735 0.920 ;
    END
END EDFKCND4

MACRO EDFKCNQD1
    CLASS CORE ;
    FOREIGN EDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.690 1.410 6.810 1.810 ;
        RECT  6.690 0.710 6.810 0.870 ;
        RECT  6.810 0.710 6.910 1.810 ;
        RECT  6.910 0.710 6.950 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 2.230 0.300 ;
        RECT  2.230 -0.300 2.450 0.340 ;
        RECT  2.450 -0.300 2.760 0.300 ;
        RECT  2.760 -0.300 2.980 0.340 ;
        RECT  2.980 -0.300 4.430 0.300 ;
        RECT  4.430 -0.300 4.650 0.480 ;
        RECT  4.650 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 2.760 2.820 ;
        RECT  2.760 2.180 2.980 2.820 ;
        RECT  2.980 2.220 4.430 2.820 ;
        RECT  4.430 1.960 4.650 2.820 ;
        RECT  4.650 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.210 0.730 5.330 1.520 ;
        RECT  5.230 0.450 5.450 0.610 ;
        RECT  5.770 0.830 6.340 0.990 ;
        RECT  1.730 1.230 1.890 1.810 ;
        RECT  1.890 1.690 4.830 1.810 ;
        RECT  4.830 1.690 4.950 2.050 ;
        RECT  4.950 1.930 5.610 2.050 ;
        RECT  5.610 1.930 5.830 2.090 ;
        RECT  5.690 0.470 5.830 0.710 ;
        RECT  5.830 1.930 7.070 2.050 ;
        RECT  5.830 0.470 7.070 0.590 ;
        RECT  7.070 0.470 7.190 2.050 ;
        RECT  6.310 1.650 6.450 1.810 ;
        RECT  6.340 0.710 6.450 0.990 ;
        RECT  6.450 0.710 6.560 1.810 ;
        RECT  6.560 0.830 6.570 1.810 ;
        RECT  6.570 1.080 6.690 1.240 ;
        RECT  5.450 0.450 5.570 1.240 ;
        RECT  5.190 1.650 5.800 1.810 ;
        RECT  5.570 1.120 5.800 1.240 ;
        RECT  5.800 1.120 5.920 1.810 ;
        RECT  5.920 1.120 6.320 1.280 ;
        RECT  5.330 1.360 5.680 1.520 ;
        RECT  4.550 1.410 4.970 1.570 ;
        RECT  4.810 0.580 4.970 0.740 ;
        RECT  4.970 0.580 5.090 1.570 ;
        RECT  3.910 0.530 4.070 1.570 ;
        RECT  4.070 0.860 4.710 0.980 ;
        RECT  4.710 0.860 4.850 1.290 ;
        RECT  1.450 0.470 3.500 0.590 ;
        RECT  3.500 0.430 3.740 0.590 ;
        RECT  3.160 0.710 3.550 0.860 ;
        RECT  3.550 0.710 3.710 1.570 ;
        RECT  1.360 1.930 2.210 2.050 ;
        RECT  2.210 1.930 2.430 2.090 ;
        RECT  2.430 1.930 3.430 2.050 ;
        RECT  3.430 1.930 3.670 2.090 ;
        RECT  2.450 0.710 2.920 0.860 ;
        RECT  2.920 0.710 3.040 1.570 ;
        RECT  3.040 1.030 3.180 1.190 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  4.390 1.100 4.550 1.570 ;
        RECT  3.830 1.410 3.910 1.570 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  3.160 1.410 3.550 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.450 1.410 2.920 1.570 ;
        RECT  0.190 1.510 0.350 1.900 ;
    END
END EDFKCNQD1

MACRO EDFKCNQD2
    CLASS CORE ;
    FOREIGN EDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.225 1.410 7.445 1.810 ;
        RECT  7.445 1.410 7.450 1.530 ;
        RECT  7.205 0.710 7.450 0.870 ;
        RECT  7.450 0.710 7.590 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 2.230 0.300 ;
        RECT  2.230 -0.300 2.450 0.340 ;
        RECT  2.450 -0.300 2.855 0.300 ;
        RECT  2.855 -0.300 3.075 0.340 ;
        RECT  3.075 -0.300 4.545 0.300 ;
        RECT  4.545 -0.300 4.765 0.480 ;
        RECT  4.765 -0.300 7.625 0.300 ;
        RECT  7.625 -0.300 7.845 0.340 ;
        RECT  7.845 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 2.855 2.820 ;
        RECT  2.855 2.180 3.075 2.820 ;
        RECT  3.075 2.220 4.545 2.820 ;
        RECT  4.545 2.040 4.765 2.820 ;
        RECT  4.765 2.220 7.625 2.820 ;
        RECT  7.625 2.180 7.845 2.820 ;
        RECT  7.845 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.085 0.580 5.205 1.570 ;
        RECT  4.025 0.530 4.185 1.570 ;
        RECT  4.185 0.860 4.825 0.980 ;
        RECT  4.825 0.860 4.965 1.290 ;
        RECT  1.450 0.470 3.595 0.590 ;
        RECT  3.595 0.430 3.835 0.590 ;
        RECT  3.255 0.710 3.645 0.860 ;
        RECT  3.645 0.710 3.805 1.570 ;
        RECT  1.360 1.930 2.210 2.050 ;
        RECT  2.210 1.930 2.430 2.090 ;
        RECT  2.430 1.930 3.525 2.050 ;
        RECT  3.525 1.930 3.765 2.090 ;
        RECT  2.545 0.710 3.015 0.860 ;
        RECT  3.015 0.710 3.135 1.570 ;
        RECT  3.135 1.030 3.275 1.190 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  4.925 0.580 5.085 0.740 ;
        RECT  4.665 1.410 5.085 1.570 ;
        RECT  5.445 1.410 5.795 1.550 ;
        RECT  6.035 1.140 6.445 1.280 ;
        RECT  5.915 1.140 6.035 1.810 ;
        RECT  5.685 1.140 5.915 1.260 ;
        RECT  5.305 1.680 5.915 1.810 ;
        RECT  5.565 0.450 5.685 1.260 ;
        RECT  6.695 1.080 7.265 1.240 ;
        RECT  6.575 0.750 6.695 1.810 ;
        RECT  6.465 0.750 6.575 1.010 ;
        RECT  6.455 1.400 6.575 1.810 ;
        RECT  7.730 0.470 7.850 2.050 ;
        RECT  5.945 0.470 7.730 0.590 ;
        RECT  5.945 1.930 7.730 2.050 ;
        RECT  5.805 0.470 5.945 0.740 ;
        RECT  5.725 1.930 5.945 2.090 ;
        RECT  5.065 1.930 5.725 2.050 ;
        RECT  4.945 1.690 5.065 2.050 ;
        RECT  1.890 1.690 4.945 1.810 ;
        RECT  5.875 0.885 6.465 1.010 ;
        RECT  5.325 0.450 5.565 0.610 ;
        RECT  5.325 0.740 5.445 1.550 ;
        RECT  4.505 1.100 4.665 1.570 ;
        RECT  3.945 1.410 4.025 1.570 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  3.255 1.410 3.645 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.545 1.410 3.015 1.570 ;
        RECT  0.190 1.510 0.350 1.900 ;
        RECT  1.730 1.230 1.890 1.810 ;
    END
END EDFKCNQD2

MACRO EDFKCNQD4
    CLASS CORE ;
    FOREIGN EDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.180 1.580 7.630 1.740 ;
        RECT  7.180 0.760 7.630 0.920 ;
        RECT  7.630 0.760 8.050 1.740 ;
        RECT  8.050 1.580 8.130 1.740 ;
        RECT  8.050 0.760 8.130 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.390 ;
        RECT  1.190 1.230 1.270 1.390 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.210 1.270 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.340 ;
        RECT  0.570 -0.300 4.445 0.300 ;
        RECT  4.445 -0.300 4.665 0.480 ;
        RECT  4.665 -0.300 6.055 0.300 ;
        RECT  6.055 -0.300 6.275 0.340 ;
        RECT  6.275 -0.300 8.290 0.300 ;
        RECT  8.290 -0.300 8.510 0.340 ;
        RECT  8.510 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.750 0.760 2.820 ;
        RECT  0.760 2.220 1.820 2.820 ;
        RECT  1.820 2.180 2.040 2.820 ;
        RECT  2.040 2.220 4.445 2.820 ;
        RECT  4.445 2.040 4.665 2.820 ;
        RECT  4.665 2.220 6.045 2.820 ;
        RECT  6.045 2.180 6.265 2.820 ;
        RECT  6.265 2.220 8.290 2.820 ;
        RECT  8.290 2.180 8.510 2.820 ;
        RECT  8.510 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.985 0.580 5.105 1.570 ;
        RECT  3.920 0.430 4.080 1.570 ;
        RECT  4.080 0.860 4.725 0.980 ;
        RECT  4.725 0.860 4.865 1.290 ;
        RECT  1.310 0.470 1.450 0.880 ;
        RECT  1.450 0.470 3.510 0.590 ;
        RECT  3.510 0.430 3.750 0.590 ;
        RECT  3.170 0.710 3.560 0.860 ;
        RECT  3.560 0.710 3.720 1.570 ;
        RECT  1.360 1.930 2.220 2.050 ;
        RECT  2.220 1.930 2.440 2.090 ;
        RECT  2.440 1.930 3.440 2.050 ;
        RECT  3.440 1.930 3.680 2.090 ;
        RECT  2.460 0.710 2.930 0.860 ;
        RECT  2.930 0.710 3.050 1.560 ;
        RECT  3.050 1.030 3.190 1.190 ;
        RECT  0.350 1.510 0.700 1.630 ;
        RECT  0.060 0.710 0.700 0.870 ;
        RECT  0.700 0.710 0.860 1.630 ;
        RECT  0.860 1.510 1.410 1.630 ;
        RECT  1.410 1.020 1.570 1.630 ;
        RECT  4.825 0.580 4.985 0.740 ;
        RECT  4.565 1.410 4.985 1.570 ;
        RECT  5.345 1.380 5.695 1.520 ;
        RECT  5.935 1.140 6.445 1.260 ;
        RECT  5.815 1.140 5.935 1.810 ;
        RECT  5.585 1.140 5.815 1.260 ;
        RECT  5.205 1.650 5.815 1.810 ;
        RECT  5.465 0.450 5.585 1.260 ;
        RECT  6.715 1.050 7.240 1.270 ;
        RECT  6.685 0.830 6.715 1.810 ;
        RECT  6.575 0.710 6.685 1.810 ;
        RECT  6.455 0.710 6.575 1.020 ;
        RECT  6.435 1.650 6.575 1.810 ;
        RECT  8.350 0.470 8.470 2.050 ;
        RECT  5.845 0.470 8.350 0.590 ;
        RECT  5.845 1.930 8.350 2.050 ;
        RECT  5.705 0.470 5.845 0.710 ;
        RECT  5.625 1.930 5.845 2.090 ;
        RECT  4.965 1.930 5.625 2.050 ;
        RECT  4.845 1.690 4.965 2.050 ;
        RECT  1.890 1.690 4.845 1.810 ;
        RECT  1.730 1.230 1.890 1.810 ;
        RECT  5.765 0.880 6.455 1.020 ;
        RECT  5.245 0.450 5.465 0.610 ;
        RECT  5.225 0.730 5.345 1.520 ;
        RECT  4.405 1.100 4.565 1.570 ;
        RECT  3.840 1.410 3.920 1.570 ;
        RECT  3.170 1.410 3.560 1.570 ;
        RECT  1.200 1.750 1.360 2.050 ;
        RECT  2.460 1.400 2.930 1.560 ;
        RECT  0.190 1.510 0.350 1.900 ;
        LAYER M1 ;
        RECT  7.180 1.580 7.415 1.740 ;
        RECT  7.180 0.760 7.415 0.920 ;
    END
END EDFKCNQD4

MACRO EDFQD1
    CLASS CORE ;
    FOREIGN EDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 0.440 7.270 1.880 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.910 0.300 ;
        RECT  1.910 -0.300 2.130 0.340 ;
        RECT  2.130 -0.300 4.440 0.300 ;
        RECT  4.440 -0.300 4.660 0.720 ;
        RECT  4.660 -0.300 6.030 0.300 ;
        RECT  6.030 -0.300 6.250 0.340 ;
        RECT  6.250 -0.300 6.680 0.300 ;
        RECT  6.680 -0.300 6.900 0.340 ;
        RECT  6.900 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 1.960 2.820 ;
        RECT  1.960 2.180 2.180 2.820 ;
        RECT  2.180 2.220 2.610 2.820 ;
        RECT  2.610 2.180 2.830 2.820 ;
        RECT  2.830 2.220 4.360 2.820 ;
        RECT  4.360 1.970 4.580 2.820 ;
        RECT  4.580 2.220 5.930 2.820 ;
        RECT  5.930 2.180 6.150 2.820 ;
        RECT  6.150 2.220 6.680 2.820 ;
        RECT  6.680 2.180 6.900 2.820 ;
        RECT  6.900 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.390 0.470 5.510 1.070 ;
        RECT  5.110 1.690 5.620 1.810 ;
        RECT  5.510 0.950 5.620 1.070 ;
        RECT  5.620 0.950 5.740 1.810 ;
        RECT  5.740 1.390 6.180 1.510 ;
        RECT  6.180 1.030 6.320 1.510 ;
        RECT  5.270 1.270 5.340 1.390 ;
        RECT  5.340 1.270 5.500 1.570 ;
        RECT  4.390 1.420 4.890 1.560 ;
        RECT  4.890 0.445 5.020 1.560 ;
        RECT  3.890 0.840 4.630 0.960 ;
        RECT  4.630 0.840 4.770 1.260 ;
        RECT  2.970 0.710 3.100 0.850 ;
        RECT  3.100 0.710 3.220 1.570 ;
        RECT  3.220 1.080 3.230 1.570 ;
        RECT  3.230 1.080 3.610 1.240 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.310 2.050 ;
        RECT  3.310 1.930 3.550 2.090 ;
        RECT  3.340 0.470 3.500 0.710 ;
        RECT  2.250 0.710 2.730 0.850 ;
        RECT  2.730 0.710 2.850 1.500 ;
        RECT  2.850 1.020 2.980 1.180 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  6.560 1.050 6.750 1.270 ;
        RECT  6.440 0.710 6.560 1.810 ;
        RECT  6.020 0.710 6.440 0.870 ;
        RECT  6.310 1.650 6.440 1.810 ;
        RECT  6.870 0.470 6.990 2.050 ;
        RECT  5.850 0.470 6.870 0.590 ;
        RECT  5.770 1.930 6.870 2.050 ;
        RECT  5.630 0.420 5.850 0.590 ;
        RECT  5.550 1.930 5.770 2.090 ;
        RECT  4.930 1.930 5.550 2.050 ;
        RECT  4.810 1.690 4.930 2.050 ;
        RECT  1.990 1.690 4.810 1.810 ;
        RECT  1.830 1.360 1.990 1.810 ;
        RECT  5.860 0.710 6.020 1.270 ;
        RECT  5.240 0.470 5.390 0.630 ;
        RECT  5.140 0.750 5.270 1.390 ;
        RECT  4.230 1.080 4.390 1.560 ;
        RECT  3.730 0.530 3.890 1.570 ;
        RECT  2.990 1.410 3.100 1.570 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.340 0.590 ;
        RECT  2.230 1.360 2.730 1.500 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFQD1

MACRO EDFQD2
    CLASS CORE ;
    FOREIGN EDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.940 1.410 7.130 1.810 ;
        RECT  6.920 0.710 7.130 0.870 ;
        RECT  7.130 0.710 7.160 1.810 ;
        RECT  7.160 0.710 7.270 1.530 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 1.910 0.300 ;
        RECT  1.910 -0.300 2.130 0.340 ;
        RECT  2.130 -0.300 2.480 0.300 ;
        RECT  2.480 -0.300 2.700 0.340 ;
        RECT  2.700 -0.300 4.360 0.300 ;
        RECT  4.360 -0.300 4.580 0.720 ;
        RECT  4.580 -0.300 7.340 0.300 ;
        RECT  7.340 -0.300 7.560 0.340 ;
        RECT  7.560 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 1.960 2.820 ;
        RECT  1.960 2.180 2.180 2.820 ;
        RECT  2.180 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.280 2.820 ;
        RECT  4.280 1.970 4.500 2.820 ;
        RECT  4.500 2.220 7.340 2.820 ;
        RECT  7.340 2.180 7.560 2.820 ;
        RECT  7.560 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.230 1.650 6.625 1.810 ;
        RECT  6.040 0.710 6.625 0.850 ;
        RECT  6.625 0.710 6.745 1.810 ;
        RECT  6.745 1.080 6.965 1.240 ;
        RECT  5.320 0.470 5.440 1.070 ;
        RECT  5.030 1.690 5.540 1.810 ;
        RECT  5.440 0.950 5.540 1.070 ;
        RECT  5.540 0.950 5.660 1.810 ;
        RECT  5.660 1.390 6.250 1.510 ;
        RECT  6.250 1.030 6.410 1.510 ;
        RECT  5.200 1.270 5.260 1.390 ;
        RECT  5.260 1.270 5.420 1.570 ;
        RECT  4.310 1.420 4.810 1.560 ;
        RECT  4.810 0.445 4.940 1.560 ;
        RECT  3.650 0.530 3.810 1.560 ;
        RECT  3.810 1.400 3.840 1.560 ;
        RECT  3.810 0.840 4.550 0.960 ;
        RECT  4.550 0.840 4.690 1.260 ;
        RECT  2.890 0.710 3.020 0.850 ;
        RECT  3.020 0.710 3.140 1.570 ;
        RECT  3.140 1.080 3.150 1.570 ;
        RECT  3.150 1.080 3.530 1.240 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.230 2.050 ;
        RECT  3.230 1.930 3.470 2.090 ;
        RECT  3.260 0.470 3.420 0.710 ;
        RECT  2.170 0.710 2.650 0.850 ;
        RECT  2.650 0.710 2.770 1.560 ;
        RECT  2.770 1.080 2.900 1.240 ;
        RECT  0.060 1.720 0.280 1.880 ;
        RECT  0.280 1.720 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  5.940 0.710 6.040 1.170 ;
        RECT  5.920 0.710 5.940 1.270 ;
        RECT  7.440 0.470 7.580 2.050 ;
        RECT  5.740 0.470 7.440 0.590 ;
        RECT  5.690 1.930 7.440 2.050 ;
        RECT  5.580 0.470 5.740 0.730 ;
        RECT  5.470 1.930 5.690 2.090 ;
        RECT  4.850 1.930 5.470 2.050 ;
        RECT  4.730 1.690 4.850 2.050 ;
        RECT  1.980 1.690 4.730 1.810 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  5.780 1.050 5.920 1.270 ;
        RECT  5.160 0.470 5.320 0.630 ;
        RECT  5.060 0.750 5.200 1.390 ;
        RECT  4.150 1.080 4.310 1.560 ;
        RECT  3.620 1.400 3.650 1.560 ;
        RECT  2.910 1.410 3.020 1.570 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.260 0.590 ;
        RECT  2.190 1.420 2.650 1.560 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  0.940 1.370 0.985 1.590 ;
    END
END EDFQD2

MACRO EDFQD4
    CLASS CORE ;
    FOREIGN EDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.190 1.600 7.630 1.760 ;
        RECT  7.220 0.710 7.630 0.870 ;
        RECT  7.630 0.710 8.050 1.760 ;
        RECT  8.050 1.600 8.140 1.760 ;
        RECT  8.050 0.710 8.170 0.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.570 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.470 ;
        RECT  0.690 -0.300 4.280 0.300 ;
        RECT  4.280 -0.300 4.500 0.720 ;
        RECT  4.500 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 2.000 0.670 2.820 ;
        RECT  0.670 2.220 4.280 2.820 ;
        RECT  4.280 1.970 4.500 2.820 ;
        RECT  4.500 2.220 6.120 2.820 ;
        RECT  6.120 2.180 6.340 2.820 ;
        RECT  6.340 2.220 8.300 2.820 ;
        RECT  8.300 2.180 8.520 2.820 ;
        RECT  8.520 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.020 0.710 3.140 1.570 ;
        RECT  3.140 1.080 3.150 1.570 ;
        RECT  3.150 1.080 3.530 1.240 ;
        RECT  1.380 1.930 1.500 2.100 ;
        RECT  1.500 1.930 3.230 2.050 ;
        RECT  3.230 1.930 3.470 2.090 ;
        RECT  3.260 0.470 3.420 0.710 ;
        RECT  2.170 0.710 2.650 0.850 ;
        RECT  2.650 0.710 2.770 1.560 ;
        RECT  2.770 1.080 2.900 1.240 ;
        RECT  0.060 1.700 0.690 1.860 ;
        RECT  0.260 0.700 0.690 0.820 ;
        RECT  0.690 0.700 0.810 1.860 ;
        RECT  0.810 1.720 1.150 1.860 ;
        RECT  1.150 1.670 1.270 1.860 ;
        RECT  1.270 1.670 1.410 1.790 ;
        RECT  1.410 1.060 1.570 1.790 ;
        RECT  0.930 0.540 0.985 0.780 ;
        RECT  0.985 0.540 1.060 1.590 ;
        RECT  1.060 0.540 1.105 1.520 ;
        RECT  2.890 0.710 3.020 0.850 ;
        RECT  4.470 0.840 4.610 1.260 ;
        RECT  3.810 0.840 4.470 0.960 ;
        RECT  3.810 1.400 3.840 1.560 ;
        RECT  3.650 0.530 3.810 1.560 ;
        RECT  3.620 1.400 3.650 1.560 ;
        RECT  4.870 1.425 4.890 1.560 ;
        RECT  4.730 0.540 4.870 1.560 ;
        RECT  4.310 1.420 4.730 1.560 ;
        RECT  4.150 1.080 4.310 1.560 ;
        RECT  6.520 1.030 6.680 1.510 ;
        RECT  5.280 1.390 6.520 1.510 ;
        RECT  5.160 0.590 5.280 1.810 ;
        RECT  5.040 0.590 5.160 0.750 ;
        RECT  7.045 1.080 7.305 1.240 ;
        RECT  6.925 0.730 7.045 1.810 ;
        RECT  6.180 0.730 6.925 0.850 ;
        RECT  6.500 1.650 6.925 1.810 ;
        RECT  6.060 0.730 6.180 1.240 ;
        RECT  8.350 0.470 8.490 2.050 ;
        RECT  5.630 0.470 8.350 0.590 ;
        RECT  5.690 1.930 8.350 2.050 ;
        RECT  5.470 1.930 5.690 2.090 ;
        RECT  5.470 0.470 5.630 0.800 ;
        RECT  4.850 1.930 5.470 2.050 ;
        RECT  4.730 1.690 4.850 2.050 ;
        RECT  1.980 1.690 4.730 1.810 ;
        RECT  5.940 1.080 6.060 1.240 ;
        RECT  5.030 1.650 5.160 1.810 ;
        RECT  2.910 1.410 3.020 1.570 ;
        RECT  1.260 1.980 1.380 2.100 ;
        RECT  1.240 0.470 3.260 0.590 ;
        RECT  2.190 1.420 2.650 1.560 ;
        RECT  0.100 0.510 0.260 0.820 ;
        RECT  1.830 1.360 1.980 1.810 ;
        RECT  0.940 1.370 0.985 1.590 ;
        LAYER M1 ;
        RECT  7.220 0.710 7.415 0.870 ;
        RECT  7.190 1.600 7.415 1.760 ;
    END
END EDFQD4

MACRO FA1D1
    CLASS CORE ;
    FOREIGN FA1D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.720 1.960 7.750 2.100 ;
        RECT  7.750 0.420 7.910 2.100 ;
        RECT  7.910 1.960 7.940 2.100 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.960 1.410 7.130 1.550 ;
        RECT  6.980 0.450 7.130 0.870 ;
        RECT  7.130 0.450 7.200 1.550 ;
        RECT  7.200 0.750 7.270 1.550 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 0.725 6.310 1.290 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.030 3.290 1.405 ;
        RECT  3.290 1.285 3.430 1.795 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.000 0.560 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 0.470 3.760 0.690 ;
        RECT  3.760 0.470 3.880 1.630 ;
        RECT  3.880 1.040 3.910 1.260 ;
        RECT  2.260 0.470 2.360 0.660 ;
        RECT  2.260 1.610 2.380 1.770 ;
        RECT  2.360 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.530 1.160 ;
        RECT  3.530 1.020 3.640 1.160 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.930 0.800 2.050 ;
        RECT  0.640 0.760 0.800 0.880 ;
        RECT  0.800 0.760 0.920 2.050 ;
        RECT  0.920 1.080 1.480 1.240 ;
        RECT  0.920 1.930 2.550 2.050 ;
        RECT  2.540 0.710 2.550 0.870 ;
        RECT  2.550 0.710 2.690 2.050 ;
        RECT  2.690 1.470 2.710 2.050 ;
        RECT  2.690 0.710 2.780 0.870 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.090 1.610 1.860 1.770 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.770 ;
        RECT  4.030 0.620 4.150 2.050 ;
        RECT  4.000 0.620 4.030 0.860 ;
        RECT  3.940 1.830 4.030 2.050 ;
        RECT  3.050 1.930 3.940 2.050 ;
        RECT  3.030 0.710 3.150 0.870 ;
        RECT  3.030 1.570 3.050 2.050 ;
        RECT  2.910 0.710 3.030 2.050 ;
        RECT  2.890 1.000 2.910 2.050 ;
        RECT  5.670 0.710 5.800 0.850 ;
        RECT  5.550 0.710 5.670 1.540 ;
        RECT  6.570 0.470 6.690 1.550 ;
        RECT  6.470 0.470 6.570 0.590 ;
        RECT  5.940 1.410 6.570 1.550 ;
        RECT  6.250 0.430 6.470 0.590 ;
        RECT  4.950 0.470 6.250 0.590 ;
        RECT  5.800 1.030 5.940 1.550 ;
        RECT  4.790 0.470 4.950 1.760 ;
        RECT  6.790 1.910 7.030 2.070 ;
        RECT  4.480 1.910 6.790 2.050 ;
        RECT  4.480 0.570 4.540 1.690 ;
        RECT  4.380 0.570 4.480 2.050 ;
        RECT  7.590 1.030 7.630 1.270 ;
        RECT  7.470 1.030 7.590 1.790 ;
        RECT  5.260 1.670 7.470 1.790 ;
        RECT  5.260 0.710 5.400 0.850 ;
        RECT  5.100 0.710 5.260 1.790 ;
        RECT  4.320 1.570 4.380 2.050 ;
        RECT  4.660 1.600 4.790 1.760 ;
        RECT  5.430 1.400 5.550 1.540 ;
        RECT  2.810 1.000 2.890 1.220 ;
        RECT  3.620 1.410 3.760 1.630 ;
        RECT  2.140 0.470 2.260 1.770 ;
        RECT  0.420 1.635 0.640 2.050 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END FA1D1

MACRO FA1D2
    CLASS CORE ;
    FOREIGN FA1D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.960 7.670 2.100 ;
        RECT  7.670 1.390 7.770 2.100 ;
        RECT  7.670 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.830 2.100 ;
        RECT  7.830 1.960 7.860 2.100 ;
        RECT  7.830 0.780 7.910 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.920 1.960 6.950 2.100 ;
        RECT  6.950 1.390 7.110 2.100 ;
        RECT  7.110 1.390 7.130 1.515 ;
        RECT  6.930 0.710 7.130 0.870 ;
        RECT  7.110 1.960 7.140 2.100 ;
        RECT  7.130 0.710 7.270 1.515 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.330 1.515 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.030 3.290 1.405 ;
        RECT  3.290 1.285 3.430 1.795 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.000 0.560 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 0.470 2.360 0.660 ;
        RECT  2.260 1.610 2.380 1.770 ;
        RECT  2.360 0.470 3.410 0.590 ;
        RECT  3.410 0.470 3.530 1.160 ;
        RECT  3.530 1.020 3.640 1.160 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.930 0.800 2.050 ;
        RECT  0.640 0.760 0.800 0.880 ;
        RECT  0.800 0.760 0.920 2.050 ;
        RECT  0.920 1.080 1.480 1.240 ;
        RECT  0.920 1.930 2.550 2.050 ;
        RECT  2.540 0.710 2.550 0.870 ;
        RECT  2.550 0.710 2.690 2.050 ;
        RECT  2.690 1.470 2.710 2.050 ;
        RECT  2.690 0.710 2.780 0.870 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.090 1.610 1.860 1.770 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.770 ;
        RECT  3.880 1.040 3.910 1.260 ;
        RECT  3.760 0.470 3.880 1.630 ;
        RECT  3.650 0.470 3.760 0.690 ;
        RECT  4.030 0.620 4.150 2.050 ;
        RECT  4.000 0.620 4.030 0.860 ;
        RECT  3.940 1.830 4.030 2.050 ;
        RECT  3.050 1.930 3.940 2.050 ;
        RECT  3.030 0.710 3.150 0.870 ;
        RECT  3.030 1.570 3.050 2.050 ;
        RECT  2.910 0.710 3.030 2.050 ;
        RECT  2.890 1.000 2.910 2.050 ;
        RECT  5.670 0.710 5.800 0.870 ;
        RECT  5.550 0.710 5.670 1.570 ;
        RECT  6.050 0.710 6.500 0.870 ;
        RECT  5.940 1.650 6.460 1.810 ;
        RECT  5.940 0.710 6.050 1.170 ;
        RECT  5.930 0.710 5.940 1.810 ;
        RECT  5.790 1.050 5.930 1.810 ;
        RECT  4.880 1.690 5.790 1.810 ;
        RECT  4.880 0.620 5.000 0.780 ;
        RECT  6.780 1.090 7.010 1.250 ;
        RECT  6.660 1.090 6.780 2.050 ;
        RECT  4.480 1.930 6.660 2.050 ;
        RECT  4.480 0.570 4.540 1.690 ;
        RECT  4.380 0.570 4.480 2.050 ;
        RECT  7.550 1.090 7.650 1.250 ;
        RECT  7.430 0.470 7.550 1.250 ;
        RECT  5.340 0.470 7.430 0.590 ;
        RECT  5.300 0.470 5.340 0.810 ;
        RECT  5.180 0.470 5.300 1.570 ;
        RECT  4.320 1.570 4.380 2.050 ;
        RECT  4.720 0.620 4.880 1.810 ;
        RECT  5.430 1.400 5.550 1.570 ;
        RECT  5.050 1.410 5.180 1.570 ;
        RECT  2.810 1.000 2.890 1.220 ;
        RECT  3.620 1.410 3.760 1.630 ;
        RECT  2.140 0.470 2.260 1.770 ;
        RECT  0.420 1.635 0.640 2.050 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END FA1D2

MACRO FA1D4
    CLASS CORE ;
    FOREIGN FA1D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.870 1.650 10.190 2.030 ;
        RECT  9.870 0.490 10.190 0.870 ;
        RECT  10.190 0.490 10.610 2.030 ;
        RECT  10.610 1.650 10.780 2.030 ;
        RECT  10.610 0.490 10.780 0.870 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.490 1.650 8.910 2.030 ;
        RECT  8.470 0.710 8.910 0.870 ;
        RECT  8.910 0.710 9.330 2.030 ;
        RECT  9.330 1.650 9.410 2.030 ;
        RECT  9.330 0.710 9.420 0.870 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.760 1.005 7.920 1.515 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.030 3.930 1.405 ;
        RECT  3.930 1.030 4.030 1.795 ;
        RECT  4.030 1.285 4.070 1.795 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.670 0.300 ;
        RECT  6.670 -0.300 6.890 0.340 ;
        RECT  6.890 -0.300 11.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.600 2.820 ;
        RECT  6.600 2.180 6.820 2.820 ;
        RECT  6.820 2.220 7.400 2.820 ;
        RECT  7.400 2.180 7.620 2.820 ;
        RECT  7.620 2.220 11.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.770 1.475 3.790 2.100 ;
        RECT  3.790 1.930 3.820 2.100 ;
        RECT  3.770 0.710 3.890 0.870 ;
        RECT  3.820 1.930 4.650 2.050 ;
        RECT  4.650 1.890 4.770 2.050 ;
        RECT  4.740 0.620 4.770 0.860 ;
        RECT  4.770 0.620 4.890 2.050 ;
        RECT  4.390 0.470 4.500 0.690 ;
        RECT  4.500 0.470 4.620 1.630 ;
        RECT  4.620 1.000 4.650 1.220 ;
        RECT  3.000 0.470 3.100 0.630 ;
        RECT  3.000 1.650 3.120 1.810 ;
        RECT  3.100 0.470 4.150 0.590 ;
        RECT  4.150 0.470 4.270 1.160 ;
        RECT  4.270 1.020 4.380 1.160 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.930 0.290 2.100 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.290 1.930 0.770 2.050 ;
        RECT  0.290 0.760 0.770 0.880 ;
        RECT  0.770 1.930 0.800 2.100 ;
        RECT  0.800 1.370 0.960 2.100 ;
        RECT  0.960 1.930 0.990 2.100 ;
        RECT  0.770 0.460 0.990 0.880 ;
        RECT  0.990 1.930 1.170 2.050 ;
        RECT  0.990 0.760 1.170 0.880 ;
        RECT  1.170 0.760 1.290 2.050 ;
        RECT  1.290 1.080 1.810 1.240 ;
        RECT  1.290 1.930 3.280 2.050 ;
        RECT  3.280 0.710 3.420 2.050 ;
        RECT  3.420 1.480 3.450 2.050 ;
        RECT  3.420 0.710 3.520 0.870 ;
        RECT  1.460 0.470 1.680 0.890 ;
        RECT  1.680 0.470 2.500 0.590 ;
        RECT  1.680 1.670 2.600 1.810 ;
        RECT  2.500 0.470 2.600 0.890 ;
        RECT  2.600 0.470 2.720 1.810 ;
        RECT  2.180 0.710 2.340 1.550 ;
        RECT  2.340 1.410 2.370 1.550 ;
        RECT  2.340 1.050 2.480 1.270 ;
        RECT  3.650 0.710 3.770 2.100 ;
        RECT  3.630 1.050 3.650 2.100 ;
        RECT  3.550 1.050 3.630 1.270 ;
        RECT  6.410 0.710 7.310 0.870 ;
        RECT  6.410 1.410 7.240 1.570 ;
        RECT  6.290 0.710 6.410 1.570 ;
        RECT  7.605 0.710 8.040 0.870 ;
        RECT  7.605 1.650 8.040 1.810 ;
        RECT  7.485 0.710 7.605 1.810 ;
        RECT  7.200 1.080 7.485 1.240 ;
        RECT  5.620 1.690 7.485 1.810 ;
        RECT  5.620 0.620 5.740 0.780 ;
        RECT  8.320 1.080 8.580 1.240 ;
        RECT  8.200 1.080 8.320 2.050 ;
        RECT  5.220 1.930 8.200 2.050 ;
        RECT  5.220 0.570 5.280 1.690 ;
        RECT  5.120 0.570 5.220 2.050 ;
        RECT  9.730 1.080 9.975 1.240 ;
        RECT  9.610 0.470 9.730 1.240 ;
        RECT  6.090 0.470 9.610 0.590 ;
        RECT  6.050 0.470 6.090 0.810 ;
        RECT  5.930 0.470 6.050 1.570 ;
        RECT  5.790 1.410 5.930 1.570 ;
        RECT  5.060 1.570 5.120 2.050 ;
        RECT  5.460 0.620 5.620 1.810 ;
        RECT  6.170 1.410 6.290 1.570 ;
        RECT  3.600 1.960 3.630 2.100 ;
        RECT  4.360 1.410 4.500 1.630 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  1.440 1.650 1.680 1.810 ;
        RECT  2.150 1.410 2.180 1.550 ;
        LAYER M1 ;
        RECT  9.870 1.650 9.975 2.030 ;
        RECT  9.870 0.490 9.975 0.870 ;
        RECT  8.490 1.650 8.695 2.030 ;
        RECT  8.470 0.710 8.695 0.870 ;
    END
END FA1D4

MACRO FCICIND1
    CLASS CORE ;
    FOREIGN FCICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.060 0.780 0.090 1.685 ;
        RECT  0.090 0.780 0.100 2.095 ;
        RECT  0.100 0.420 0.180 2.095 ;
        RECT  0.180 0.420 0.250 0.900 ;
        RECT  0.180 1.565 0.260 2.095 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.565 0.550 2.075 ;
        RECT  0.550 1.565 0.615 1.685 ;
        RECT  0.615 1.065 0.755 1.685 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.950 1.860 1.515 ;
        RECT  1.860 0.950 2.650 1.070 ;
        RECT  2.650 0.950 2.810 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.520 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.890 0.300 ;
        RECT  1.890 -0.300 2.110 0.560 ;
        RECT  2.110 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.580 0.470 3.230 0.590 ;
        RECT  3.230 0.470 3.450 0.890 ;
        RECT  2.600 1.930 3.230 2.050 ;
        RECT  3.230 1.630 3.450 2.050 ;
        RECT  0.375 0.480 0.495 1.285 ;
        RECT  0.495 0.480 1.130 0.600 ;
        RECT  1.130 0.450 1.135 1.790 ;
        RECT  1.135 0.450 1.250 1.810 ;
        RECT  1.250 0.450 1.355 0.870 ;
        RECT  1.250 1.650 1.375 1.810 ;
        RECT  2.740 1.635 2.970 1.795 ;
        RECT  1.355 0.710 2.970 0.830 ;
        RECT  2.970 0.710 3.110 1.795 ;
        RECT  0.805 0.720 0.890 0.940 ;
        RECT  0.890 0.720 1.010 2.050 ;
        RECT  1.010 1.930 2.020 2.050 ;
        RECT  2.020 1.190 2.180 2.050 ;
        RECT  2.340 0.450 2.580 0.590 ;
        RECT  2.380 1.630 2.600 2.050 ;
        RECT  0.300 1.065 0.375 1.285 ;
        RECT  0.805 1.830 0.890 2.050 ;
    END
END FCICIND1

MACRO FCICIND2
    CLASS CORE ;
    FOREIGN FCICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.800 0.550 1.515 ;
        RECT  0.560 1.940 0.580 2.100 ;
        RECT  0.550 1.390 0.580 1.515 ;
        RECT  0.550 0.800 0.590 0.920 ;
        RECT  0.590 0.420 0.740 0.920 ;
        RECT  0.580 1.390 0.750 2.100 ;
        RECT  0.750 1.940 0.780 2.100 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.565 1.105 2.075 ;
        RECT  1.105 1.065 1.190 2.075 ;
        RECT  1.190 1.065 1.245 1.685 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.190 0.950 2.350 1.390 ;
        RECT  2.350 0.950 2.970 1.070 ;
        RECT  2.970 0.950 3.130 1.390 ;
        RECT  3.130 1.005 3.430 1.235 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 2.380 0.300 ;
        RECT  2.380 -0.300 2.600 0.560 ;
        RECT  2.600 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 2.380 2.820 ;
        RECT  2.380 2.180 2.600 2.820 ;
        RECT  2.600 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.510 1.190 2.670 1.795 ;
        RECT  2.340 1.675 2.510 1.795 ;
        RECT  2.220 1.675 2.340 2.050 ;
        RECT  1.500 1.930 2.220 2.050 ;
        RECT  1.380 0.720 1.500 2.050 ;
        RECT  1.295 0.720 1.380 0.940 ;
        RECT  3.550 0.710 3.690 1.795 ;
        RECT  2.070 0.710 3.550 0.830 ;
        RECT  3.230 1.635 3.550 1.795 ;
        RECT  1.950 0.710 2.070 1.810 ;
        RECT  1.845 0.710 1.950 0.850 ;
        RECT  1.620 1.650 1.950 1.810 ;
        RECT  1.620 0.450 1.845 0.850 ;
        RECT  0.985 0.480 1.620 0.600 ;
        RECT  0.865 0.480 0.985 1.270 ;
        RECT  3.090 1.930 3.870 2.050 ;
        RECT  3.070 0.470 3.870 0.590 ;
        RECT  2.870 1.630 3.090 2.050 ;
        RECT  0.790 1.050 0.865 1.270 ;
        RECT  1.315 1.830 1.380 2.050 ;
        RECT  2.830 0.450 3.070 0.590 ;
    END
END FCICIND2

MACRO FCICOND1
    CLASS CORE ;
    FOREIGN FCICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.450 0.610 2.070 ;
        RECT  0.610 1.650 0.715 2.070 ;
        RECT  0.610 0.450 0.715 0.870 ;
        RECT  2.100 1.635 2.330 1.795 ;
        RECT  0.715 0.710 2.330 0.830 ;
        RECT  2.330 0.710 2.470 1.795 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.190 1.540 1.795 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.950 1.220 1.795 ;
        RECT  1.220 0.950 2.010 1.070 ;
        RECT  2.010 0.950 2.170 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.880 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.560 ;
        RECT  1.470 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.590 1.630 2.810 2.050 ;
        RECT  1.960 1.930 2.590 2.050 ;
        RECT  2.590 0.470 2.810 0.890 ;
        RECT  1.940 0.470 2.590 0.590 ;
        RECT  1.700 0.450 1.940 0.590 ;
        RECT  1.740 1.630 1.960 2.050 ;
    END
END FCICOND1

MACRO FCICOND2
    CLASS CORE ;
    FOREIGN FCICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.780 0.230 1.795 ;
        RECT  0.230 1.635 0.560 1.795 ;
        RECT  0.230 0.780 0.560 0.900 ;
        RECT  0.560 1.635 0.780 2.055 ;
        RECT  0.560 0.480 0.780 0.900 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.190 2.790 1.795 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.950 2.470 1.515 ;
        RECT  2.470 0.950 3.125 1.070 ;
        RECT  3.125 0.950 3.285 1.390 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.855 1.150 2.010 1.370 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 2.365 0.300 ;
        RECT  2.365 -0.300 2.585 0.560 ;
        RECT  2.585 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 2.365 2.820 ;
        RECT  2.365 2.180 2.585 2.820 ;
        RECT  2.585 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.330 0.720 1.450 2.075 ;
        RECT  1.300 0.720 1.330 0.940 ;
        RECT  1.280 1.395 1.330 2.075 ;
        RECT  0.910 1.395 1.280 1.515 ;
        RECT  0.770 1.055 0.910 1.515 ;
        RECT  3.445 0.710 3.585 1.775 ;
        RECT  1.830 0.710 3.445 0.830 ;
        RECT  3.215 1.615 3.445 1.775 ;
        RECT  1.725 0.450 1.830 0.870 ;
        RECT  1.725 1.650 1.830 2.070 ;
        RECT  1.605 0.450 1.725 2.070 ;
        RECT  1.180 0.470 1.605 0.590 ;
        RECT  1.180 1.055 1.210 1.275 ;
        RECT  3.705 1.630 3.925 2.050 ;
        RECT  3.705 0.470 3.925 0.890 ;
        RECT  3.055 0.470 3.705 0.590 ;
        RECT  2.815 0.450 3.055 0.590 ;
        RECT  2.835 1.910 3.705 2.050 ;
        RECT  1.060 0.470 1.180 1.275 ;
        RECT  0.490 1.055 0.770 1.275 ;
    END
END FCICOND2

MACRO FCSICIND1
    CLASS CORE ;
    FOREIGN FCSICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.890 1.390 14.050 1.890 ;
        RECT  13.890 0.420 14.050 0.900 ;
        RECT  14.050 1.390 14.170 1.515 ;
        RECT  14.050 0.780 14.170 0.900 ;
        RECT  14.170 0.780 14.310 1.515 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  13.260 1.060 13.320 1.280 ;
        RECT  13.320 0.835 13.440 1.280 ;
        RECT  13.440 0.835 13.530 0.955 ;
        RECT  13.530 0.445 13.670 0.955 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 0.720 7.770 1.150 ;
        RECT  7.770 0.720 7.870 1.810 ;
        RECT  7.870 1.015 7.910 1.810 ;
        RECT  7.910 1.670 8.075 1.810 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.125 1.670 7.130 1.810 ;
        RECT  7.130 1.565 7.225 1.810 ;
        RECT  7.225 1.005 7.310 1.810 ;
        RECT  7.310 0.720 7.345 1.810 ;
        RECT  7.345 0.720 7.530 1.150 ;
        RECT  7.345 1.565 7.590 1.810 ;
        END
    END CO0
    PIN CIN1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.650 1.005 11.160 1.235 ;
        END
    END CIN1
    PIN CIN0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 0.725 4.070 1.235 ;
        RECT  4.070 1.070 4.300 1.235 ;
        END
    END CIN0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.710 0.300 ;
        RECT  6.710 -0.300 6.830 0.540 ;
        RECT  6.830 -0.300 8.295 0.300 ;
        RECT  8.295 -0.300 8.415 0.540 ;
        RECT  8.415 -0.300 14.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 14.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.800 0.470 4.920 1.570 ;
        RECT  4.920 1.430 5.080 1.570 ;
        RECT  4.920 0.470 6.470 0.590 ;
        RECT  6.470 0.470 6.590 0.790 ;
        RECT  6.590 0.670 6.950 0.790 ;
        RECT  6.950 0.470 7.070 0.790 ;
        RECT  7.070 0.470 8.055 0.590 ;
        RECT  8.055 0.470 8.175 0.790 ;
        RECT  8.175 0.670 8.535 0.790 ;
        RECT  8.535 0.470 8.655 0.790 ;
        RECT  8.655 0.470 12.620 0.590 ;
        RECT  12.620 0.470 12.710 1.810 ;
        RECT  12.710 0.420 12.740 1.810 ;
        RECT  12.740 1.640 12.900 1.810 ;
        RECT  12.740 0.420 12.950 0.590 ;
        RECT  10.390 1.930 11.880 2.050 ;
        RECT  11.880 1.830 11.920 2.050 ;
        RECT  11.920 0.710 12.040 2.050 ;
        RECT  12.040 0.710 12.090 0.930 ;
        RECT  9.870 0.710 9.990 1.810 ;
        RECT  9.990 0.710 10.130 0.930 ;
        RECT  9.990 1.690 11.500 1.810 ;
        RECT  11.500 1.670 11.640 1.810 ;
        RECT  11.610 0.710 11.640 0.930 ;
        RECT  11.640 0.710 11.760 1.810 ;
        RECT  10.790 0.715 11.280 0.875 ;
        RECT  11.280 0.715 11.400 1.570 ;
        RECT  11.400 1.040 11.520 1.260 ;
        RECT  10.260 0.710 10.380 1.570 ;
        RECT  10.380 0.710 10.510 0.940 ;
        RECT  8.245 1.260 8.310 1.810 ;
        RECT  8.310 1.380 8.365 1.810 ;
        RECT  8.365 1.690 9.370 1.810 ;
        RECT  9.370 1.590 9.410 1.810 ;
        RECT  9.410 1.120 9.530 1.810 ;
        RECT  9.530 1.120 9.540 1.260 ;
        RECT  9.540 0.710 9.660 1.260 ;
        RECT  9.660 0.710 9.750 0.940 ;
        RECT  9.090 0.730 9.220 1.570 ;
        RECT  9.220 0.730 9.420 0.900 ;
        RECT  2.860 0.710 2.980 2.050 ;
        RECT  2.980 1.630 3.080 2.050 ;
        RECT  2.980 0.710 3.130 0.870 ;
        RECT  3.080 1.930 6.020 2.050 ;
        RECT  6.020 1.930 6.240 2.070 ;
        RECT  6.240 1.930 8.940 2.050 ;
        RECT  8.940 1.930 9.180 2.070 ;
        RECT  8.700 1.030 8.810 1.570 ;
        RECT  8.810 0.720 8.820 1.570 ;
        RECT  8.820 0.720 8.970 1.250 ;
        RECT  5.455 0.710 5.575 1.260 ;
        RECT  5.575 1.120 5.605 1.260 ;
        RECT  5.605 1.120 5.725 1.810 ;
        RECT  5.725 1.630 5.840 1.810 ;
        RECT  5.840 1.690 6.800 1.810 ;
        RECT  6.800 1.280 6.920 1.810 ;
        RECT  6.920 1.280 7.020 1.500 ;
        RECT  6.350 1.030 6.470 1.570 ;
        RECT  6.470 1.430 6.600 1.570 ;
        RECT  5.950 0.730 6.080 1.570 ;
        RECT  6.080 1.430 6.220 1.570 ;
        RECT  3.500 0.740 3.780 0.900 ;
        RECT  5.040 0.710 5.190 1.260 ;
        RECT  3.500 1.690 5.210 1.810 ;
        RECT  5.190 1.120 5.210 1.260 ;
        RECT  5.210 1.120 5.330 1.810 ;
        RECT  5.330 1.400 5.460 1.620 ;
        RECT  2.260 1.590 2.360 1.750 ;
        RECT  2.260 0.470 2.360 0.630 ;
        RECT  2.360 0.470 4.460 0.590 ;
        RECT  4.460 0.420 4.680 0.590 ;
        RECT  3.810 1.450 4.340 1.570 ;
        RECT  4.340 1.430 4.430 1.570 ;
        RECT  4.270 0.720 4.430 0.940 ;
        RECT  4.430 0.720 4.550 1.570 ;
        RECT  4.550 1.430 4.560 1.570 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.895 0.830 2.015 ;
        RECT  0.640 0.760 0.830 0.880 ;
        RECT  0.830 0.760 0.950 2.015 ;
        RECT  0.950 1.090 1.180 1.250 ;
        RECT  0.950 1.895 2.490 2.015 ;
        RECT  2.490 0.710 2.630 2.015 ;
        RECT  2.630 1.560 2.710 1.780 ;
        RECT  2.630 0.710 2.730 0.930 ;
        RECT  1.110 0.470 1.300 0.890 ;
        RECT  1.300 0.470 1.330 1.775 ;
        RECT  1.330 0.765 1.420 1.775 ;
        RECT  1.420 0.765 1.760 0.885 ;
        RECT  1.760 0.470 1.980 0.885 ;
        RECT  1.420 1.635 2.000 1.775 ;
        RECT  4.780 0.720 4.800 1.570 ;
        RECT  13.140 1.400 13.260 1.590 ;
        RECT  13.140 0.720 13.200 0.940 ;
        RECT  13.020 0.720 13.140 1.590 ;
        RECT  12.990 0.720 13.020 1.250 ;
        RECT  13.590 1.090 13.750 2.050 ;
        RECT  12.490 1.930 13.590 2.050 ;
        RECT  12.330 0.710 12.490 2.050 ;
        RECT  12.880 1.030 12.990 1.250 ;
        RECT  12.270 1.830 12.330 2.050 ;
        RECT  4.670 0.720 4.780 0.940 ;
        RECT  10.150 1.930 10.390 2.070 ;
        RECT  9.750 1.470 9.870 1.690 ;
        RECT  10.650 1.430 11.280 1.570 ;
        RECT  10.140 1.430 10.260 1.570 ;
        RECT  8.140 1.260 8.245 1.500 ;
        RECT  8.950 1.430 9.090 1.570 ;
        RECT  2.750 1.050 2.860 1.270 ;
        RECT  8.580 1.430 8.700 1.570 ;
        RECT  5.410 0.710 5.455 0.930 ;
        RECT  6.210 0.720 6.350 1.250 ;
        RECT  5.740 0.730 5.950 0.910 ;
        RECT  3.380 0.740 3.500 1.810 ;
        RECT  2.140 0.470 2.260 1.750 ;
        RECT  3.650 1.060 3.810 1.570 ;
        RECT  0.420 1.595 0.640 2.015 ;
        RECT  1.090 1.615 1.300 1.775 ;
    END
END FCSICIND1

MACRO FCSICIND2
    CLASS CORE ;
    FOREIGN FCSICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.220 1.950 15.250 2.090 ;
        RECT  15.250 1.380 15.410 2.090 ;
        RECT  15.250 0.440 15.410 0.940 ;
        RECT  15.410 1.950 15.440 2.090 ;
        RECT  15.410 1.380 15.450 1.540 ;
        RECT  15.410 0.820 15.450 0.940 ;
        RECT  15.450 0.820 15.590 1.540 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.620 1.060 14.680 1.280 ;
        RECT  14.680 0.835 14.800 1.280 ;
        RECT  14.800 0.835 14.810 0.955 ;
        RECT  14.810 0.445 14.950 0.955 ;
        END
    END CS
    PIN CO1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.485 1.650 8.730 1.810 ;
        RECT  8.700 0.720 8.730 1.150 ;
        RECT  8.730 0.720 8.870 1.810 ;
        RECT  8.870 0.720 8.930 1.150 ;
        RECT  8.870 1.650 9.435 1.810 ;
        END
    END CO1
    PIN CO0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.105 1.650 7.450 1.810 ;
        RECT  7.450 1.030 7.590 1.810 ;
        RECT  7.590 1.030 7.620 1.150 ;
        RECT  7.620 0.720 7.840 1.150 ;
        RECT  7.590 1.650 8.055 1.810 ;
        END
    END CO0
    PIN CIN1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.930 1.005 12.500 1.235 ;
        END
    END CIN1
    PIN CIN0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 0.725 4.070 1.235 ;
        RECT  4.070 1.070 4.300 1.235 ;
        END
    END CIN0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.650 1.045 1.690 1.205 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.710 0.300 ;
        RECT  6.710 -0.300 6.830 0.540 ;
        RECT  6.830 -0.300 8.210 0.300 ;
        RECT  8.210 -0.300 8.330 0.540 ;
        RECT  8.330 -0.300 9.655 0.300 ;
        RECT  9.655 -0.300 9.775 0.540 ;
        RECT  9.775 -0.300 14.800 0.300 ;
        RECT  14.800 -0.300 15.020 0.325 ;
        RECT  15.020 -0.300 15.635 0.300 ;
        RECT  15.635 -0.300 15.855 0.340 ;
        RECT  15.855 -0.300 16.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 14.820 2.820 ;
        RECT  14.820 2.180 15.040 2.820 ;
        RECT  15.040 2.220 15.635 2.820 ;
        RECT  15.635 2.180 15.855 2.820 ;
        RECT  15.855 2.220 16.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.605 1.310 9.725 1.810 ;
        RECT  9.725 1.690 10.730 1.810 ;
        RECT  11.740 0.710 11.940 0.875 ;
        RECT  11.620 0.710 11.740 1.570 ;
        RECT  12.755 1.040 12.880 1.260 ;
        RECT  10.730 1.120 10.890 1.810 ;
        RECT  10.890 1.120 10.900 1.260 ;
        RECT  10.900 0.710 11.020 1.260 ;
        RECT  12.635 0.715 12.755 1.570 ;
        RECT  12.150 0.715 12.635 0.875 ;
        RECT  13.000 0.710 13.120 1.810 ;
        RECT  11.020 0.710 11.110 0.940 ;
        RECT  10.450 0.730 10.580 1.570 ;
        RECT  10.580 0.730 10.780 0.900 ;
        RECT  12.970 0.710 13.000 0.930 ;
        RECT  12.860 1.670 13.000 1.810 ;
        RECT  11.350 1.690 12.860 1.810 ;
        RECT  2.860 0.710 2.980 2.050 ;
        RECT  2.980 1.630 3.080 2.050 ;
        RECT  11.350 0.710 11.490 0.930 ;
        RECT  11.230 0.710 11.350 1.810 ;
        RECT  13.410 0.710 13.450 0.930 ;
        RECT  2.980 0.710 3.130 0.870 ;
        RECT  3.080 1.930 6.020 2.050 ;
        RECT  6.020 1.930 6.240 2.070 ;
        RECT  13.290 0.710 13.410 2.050 ;
        RECT  13.240 1.830 13.290 2.050 ;
        RECT  11.750 1.930 13.240 2.050 ;
        RECT  6.240 1.930 10.300 2.050 ;
        RECT  10.300 1.930 10.540 2.070 ;
        RECT  10.060 1.030 10.170 1.570 ;
        RECT  14.100 0.420 14.310 0.590 ;
        RECT  14.100 1.640 14.260 1.810 ;
        RECT  14.070 0.420 14.100 1.810 ;
        RECT  10.170 0.720 10.180 1.570 ;
        RECT  10.180 0.720 10.330 1.250 ;
        RECT  5.455 0.710 5.575 1.260 ;
        RECT  13.980 0.470 14.070 1.810 ;
        RECT  10.015 0.470 13.980 0.590 ;
        RECT  9.895 0.470 10.015 0.790 ;
        RECT  5.575 1.120 5.605 1.260 ;
        RECT  5.605 1.120 5.725 1.810 ;
        RECT  5.725 1.630 5.840 1.810 ;
        RECT  9.535 0.670 9.895 0.790 ;
        RECT  9.415 0.470 9.535 0.790 ;
        RECT  8.580 0.470 9.415 0.590 ;
        RECT  5.840 1.690 6.800 1.810 ;
        RECT  6.800 1.310 6.920 1.810 ;
        RECT  6.920 1.310 7.235 1.470 ;
        RECT  8.460 0.470 8.580 0.790 ;
        RECT  8.080 0.670 8.460 0.790 ;
        RECT  7.960 0.470 8.080 0.790 ;
        RECT  6.350 1.030 6.470 1.570 ;
        RECT  6.470 1.430 6.600 1.570 ;
        RECT  5.950 0.730 6.080 1.570 ;
        RECT  7.070 0.470 7.960 0.590 ;
        RECT  6.950 0.470 7.070 0.790 ;
        RECT  6.590 0.670 6.950 0.790 ;
        RECT  6.080 1.430 6.220 1.570 ;
        RECT  3.500 0.740 3.780 0.900 ;
        RECT  5.040 0.710 5.190 1.260 ;
        RECT  6.470 0.470 6.590 0.790 ;
        RECT  4.920 0.470 6.470 0.590 ;
        RECT  4.920 1.430 5.080 1.570 ;
        RECT  3.500 1.690 5.210 1.810 ;
        RECT  5.190 1.120 5.210 1.260 ;
        RECT  5.210 1.120 5.330 1.810 ;
        RECT  4.800 0.470 4.920 1.570 ;
        RECT  4.780 0.720 4.800 1.570 ;
        RECT  14.500 1.400 14.620 1.590 ;
        RECT  5.330 1.400 5.460 1.620 ;
        RECT  2.260 1.590 2.360 1.750 ;
        RECT  2.260 0.470 2.360 0.630 ;
        RECT  14.500 0.700 14.560 0.940 ;
        RECT  14.380 0.700 14.500 1.590 ;
        RECT  14.940 1.090 15.100 2.050 ;
        RECT  2.360 0.470 4.460 0.590 ;
        RECT  4.460 0.420 4.680 0.590 ;
        RECT  3.810 1.450 4.340 1.570 ;
        RECT  13.850 1.930 14.940 2.050 ;
        RECT  13.690 0.710 13.850 2.050 ;
        RECT  4.340 1.430 4.430 1.570 ;
        RECT  4.270 0.720 4.430 0.940 ;
        RECT  4.430 0.720 4.550 1.570 ;
        RECT  4.550 1.430 4.560 1.570 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.895 0.830 2.015 ;
        RECT  0.640 0.760 0.830 0.880 ;
        RECT  0.830 0.760 0.950 2.015 ;
        RECT  0.950 1.090 1.180 1.250 ;
        RECT  0.950 1.895 2.490 2.015 ;
        RECT  2.490 0.710 2.630 2.015 ;
        RECT  2.630 1.560 2.710 1.780 ;
        RECT  2.630 0.710 2.730 0.930 ;
        RECT  1.110 0.470 1.300 0.890 ;
        RECT  1.300 0.470 1.330 1.775 ;
        RECT  1.330 0.765 1.420 1.775 ;
        RECT  1.420 0.765 1.760 0.885 ;
        RECT  1.760 0.470 1.980 0.885 ;
        RECT  1.420 1.635 2.000 1.775 ;
        RECT  14.240 1.030 14.380 1.250 ;
        RECT  13.630 1.830 13.690 2.050 ;
        RECT  4.670 0.720 4.780 0.940 ;
        RECT  11.510 1.930 11.750 2.070 ;
        RECT  11.110 1.500 11.230 1.720 ;
        RECT  11.950 1.430 12.635 1.570 ;
        RECT  11.500 1.430 11.620 1.570 ;
        RECT  9.305 1.310 9.605 1.470 ;
        RECT  10.310 1.430 10.450 1.570 ;
        RECT  2.750 1.050 2.860 1.270 ;
        RECT  9.940 1.430 10.060 1.570 ;
        RECT  5.410 0.710 5.455 0.940 ;
        RECT  6.210 0.720 6.350 1.250 ;
        RECT  5.740 0.730 5.950 0.910 ;
        RECT  3.380 0.740 3.500 1.810 ;
        RECT  2.140 0.470 2.260 1.750 ;
        RECT  3.650 1.060 3.810 1.570 ;
        RECT  0.420 1.595 0.640 2.015 ;
        RECT  1.090 1.615 1.300 1.775 ;
    END
END FCSICIND2

MACRO FCSICOND1
    CLASS CORE ;
    FOREIGN FCSICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  15.230 1.565 15.390 2.095 ;
        RECT  15.230 0.420 15.390 0.900 ;
        RECT  15.390 1.565 15.450 1.685 ;
        RECT  15.390 0.780 15.450 0.900 ;
        RECT  15.450 0.780 15.590 1.685 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.545 1.060 14.595 1.300 ;
        RECT  14.595 0.835 14.715 1.300 ;
        RECT  14.715 0.835 14.810 0.955 ;
        RECT  14.810 0.445 14.950 0.955 ;
        END
    END CS
    PIN CON1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.410 0.915 8.550 1.810 ;
        RECT  8.550 1.670 8.820 1.810 ;
        RECT  8.550 0.915 8.995 1.075 ;
        END
    END CON1
    PIN CON0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.830 1.670 8.090 1.810 ;
        RECT  7.630 0.915 8.090 1.075 ;
        RECT  8.090 0.915 8.230 1.810 ;
        END
    END CON0
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.630 1.090 12.890 1.310 ;
        RECT  12.890 1.005 13.030 1.515 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.750 1.515 ;
        RECT  3.750 1.080 3.960 1.300 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.060 3.290 1.280 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.840 0.300 ;
        RECT  6.840 -0.300 6.960 0.520 ;
        RECT  6.960 -0.300 8.250 0.300 ;
        RECT  8.250 -0.300 8.370 0.520 ;
        RECT  8.370 -0.300 9.650 0.300 ;
        RECT  9.650 -0.300 9.770 0.520 ;
        RECT  9.770 -0.300 14.770 0.300 ;
        RECT  14.770 -0.300 14.990 0.325 ;
        RECT  14.990 -0.300 15.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 14.785 2.820 ;
        RECT  14.785 2.180 15.005 2.820 ;
        RECT  15.005 2.220 15.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.010 0.470 13.940 0.590 ;
        RECT  13.940 0.470 14.060 1.810 ;
        RECT  14.060 1.590 14.180 1.810 ;
        RECT  14.060 0.420 14.280 0.590 ;
        RECT  11.740 1.930 13.210 2.050 ;
        RECT  13.210 0.710 13.380 2.050 ;
        RECT  13.380 0.710 13.400 0.930 ;
        RECT  11.180 1.120 11.200 1.690 ;
        RECT  11.200 1.120 11.320 1.810 ;
        RECT  11.320 1.120 11.340 1.260 ;
        RECT  11.340 0.710 11.500 1.260 ;
        RECT  11.320 1.690 12.300 1.810 ;
        RECT  12.300 0.760 12.460 1.810 ;
        RECT  12.460 0.760 12.860 0.880 ;
        RECT  12.460 1.670 13.070 1.810 ;
        RECT  12.860 0.740 13.080 0.880 ;
        RECT  11.680 0.740 11.820 1.570 ;
        RECT  11.820 0.740 11.930 0.900 ;
        RECT  9.590 1.080 9.710 1.810 ;
        RECT  9.710 1.690 10.720 1.810 ;
        RECT  10.720 1.590 10.790 1.810 ;
        RECT  10.790 1.120 10.910 1.810 ;
        RECT  10.910 1.120 10.940 1.260 ;
        RECT  10.940 0.710 11.060 1.260 ;
        RECT  11.060 0.710 11.120 0.940 ;
        RECT  10.470 0.730 10.600 1.570 ;
        RECT  10.600 0.730 10.790 0.910 ;
        RECT  2.890 1.050 2.900 2.050 ;
        RECT  2.900 0.760 3.030 2.050 ;
        RECT  3.030 1.470 3.050 2.050 ;
        RECT  3.030 0.760 3.140 0.920 ;
        RECT  3.050 1.930 6.150 2.050 ;
        RECT  6.150 1.930 6.370 2.070 ;
        RECT  6.370 1.930 10.290 2.050 ;
        RECT  10.290 1.930 10.530 2.070 ;
        RECT  10.060 1.090 10.130 1.570 ;
        RECT  10.130 0.720 10.180 1.570 ;
        RECT  10.180 0.720 10.270 1.210 ;
        RECT  10.270 0.990 10.350 1.210 ;
        RECT  9.150 0.720 9.290 1.810 ;
        RECT  9.290 1.670 9.460 1.810 ;
        RECT  7.320 0.720 7.440 1.810 ;
        RECT  7.440 0.720 7.460 1.505 ;
        RECT  7.460 1.345 7.720 1.505 ;
        RECT  5.600 0.710 5.720 1.260 ;
        RECT  5.720 1.120 5.780 1.260 ;
        RECT  5.780 1.120 5.920 1.810 ;
        RECT  5.920 1.690 6.870 1.810 ;
        RECT  6.870 1.180 6.980 1.810 ;
        RECT  6.980 1.060 6.990 1.810 ;
        RECT  6.990 1.060 7.150 1.300 ;
        RECT  6.340 0.720 6.480 1.250 ;
        RECT  6.480 1.130 6.600 1.570 ;
        RECT  6.600 1.430 6.730 1.570 ;
        RECT  6.040 0.740 6.170 1.570 ;
        RECT  6.170 1.430 6.350 1.570 ;
        RECT  3.770 1.690 4.080 1.810 ;
        RECT  3.530 0.710 4.080 0.870 ;
        RECT  4.080 0.710 4.200 1.810 ;
        RECT  4.200 1.050 4.340 1.210 ;
        RECT  5.170 0.710 5.320 1.260 ;
        RECT  4.200 1.690 5.340 1.810 ;
        RECT  5.320 1.120 5.340 1.260 ;
        RECT  5.340 1.120 5.460 1.810 ;
        RECT  5.460 1.120 5.480 1.680 ;
        RECT  5.480 1.520 5.610 1.680 ;
        RECT  2.260 0.470 2.360 0.630 ;
        RECT  2.260 1.590 2.380 1.750 ;
        RECT  2.360 0.470 4.590 0.590 ;
        RECT  4.590 0.420 4.810 0.590 ;
        RECT  4.320 0.760 4.505 0.920 ;
        RECT  4.505 0.760 4.625 1.560 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.895 0.850 2.015 ;
        RECT  0.640 0.760 0.850 0.880 ;
        RECT  0.850 0.760 0.990 2.015 ;
        RECT  0.990 1.090 1.460 1.250 ;
        RECT  0.990 1.895 2.550 2.015 ;
        RECT  2.540 0.710 2.550 0.830 ;
        RECT  2.550 0.710 2.690 2.015 ;
        RECT  2.690 1.470 2.710 2.015 ;
        RECT  2.690 0.710 2.780 0.850 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.110 1.570 1.860 1.730 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.730 ;
        RECT  9.890 0.470 10.010 0.760 ;
        RECT  9.530 0.640 9.890 0.760 ;
        RECT  9.410 0.470 9.530 0.760 ;
        RECT  8.610 0.470 9.410 0.590 ;
        RECT  8.490 0.470 8.610 0.760 ;
        RECT  8.130 0.640 8.490 0.760 ;
        RECT  8.010 0.470 8.130 0.760 ;
        RECT  7.200 0.470 8.010 0.590 ;
        RECT  7.080 0.470 7.200 0.760 ;
        RECT  6.720 0.640 7.080 0.760 ;
        RECT  6.600 0.470 6.720 0.760 ;
        RECT  5.050 0.470 6.600 0.590 ;
        RECT  5.050 1.430 5.210 1.570 ;
        RECT  4.930 0.470 5.050 1.570 ;
        RECT  4.910 0.710 4.930 1.570 ;
        RECT  14.420 1.430 14.600 1.590 ;
        RECT  14.420 0.720 14.475 0.940 ;
        RECT  14.300 0.720 14.420 1.590 ;
        RECT  15.090 1.090 15.140 1.310 ;
        RECT  14.970 1.090 15.090 1.870 ;
        RECT  14.535 1.750 14.970 1.870 ;
        RECT  14.415 1.750 14.535 2.050 ;
        RECT  13.820 1.930 14.415 2.050 ;
        RECT  13.740 1.890 13.820 2.050 ;
        RECT  13.740 0.710 13.810 0.940 ;
        RECT  14.180 1.030 14.300 1.250 ;
        RECT  4.750 0.710 4.910 0.930 ;
        RECT  11.500 1.930 11.740 2.070 ;
        RECT  11.050 1.530 11.180 1.690 ;
        RECT  11.450 1.430 11.680 1.570 ;
        RECT  9.510 1.080 9.590 1.300 ;
        RECT  10.310 1.430 10.470 1.570 ;
        RECT  2.810 1.050 2.890 1.270 ;
        RECT  9.930 1.430 10.060 1.570 ;
        RECT  8.830 1.345 9.150 1.505 ;
        RECT  7.170 1.670 7.320 1.810 ;
        RECT  5.540 0.710 5.600 0.940 ;
        RECT  6.290 1.030 6.340 1.250 ;
        RECT  5.870 0.740 6.040 0.900 ;
        RECT  3.530 1.670 3.770 1.810 ;
        RECT  2.140 0.470 2.260 1.750 ;
        RECT  4.350 1.400 4.505 1.560 ;
        RECT  0.420 1.595 0.640 2.015 ;
        RECT  13.600 0.710 13.740 2.050 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END FCSICOND1

MACRO FCSICOND2
    CLASS CORE ;
    FOREIGN FCSICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  16.500 1.950 16.530 2.090 ;
        RECT  16.530 1.380 16.690 2.090 ;
        RECT  16.530 0.440 16.690 0.940 ;
        RECT  16.690 1.950 16.720 2.090 ;
        RECT  16.690 1.380 16.730 1.540 ;
        RECT  16.690 0.790 16.730 0.940 ;
        RECT  16.730 0.790 16.870 1.540 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  15.925 1.060 15.975 1.300 ;
        RECT  15.975 0.835 16.090 1.300 ;
        RECT  16.090 0.445 16.095 1.300 ;
        RECT  16.095 0.445 16.230 0.955 ;
        END
    END CS
    PIN CON1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.250 1.670 9.370 1.810 ;
        RECT  9.120 0.915 9.370 1.075 ;
        RECT  9.370 0.915 9.510 1.810 ;
        RECT  9.510 1.670 10.240 1.810 ;
        RECT  9.510 0.915 10.415 1.075 ;
        END
    END CON1
    PIN CON0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.830 1.670 8.410 1.810 ;
        RECT  7.630 0.915 8.410 1.075 ;
        RECT  8.410 0.915 8.550 1.810 ;
        RECT  8.550 1.670 8.800 1.810 ;
        RECT  8.550 0.915 8.980 1.075 ;
        END
    END CON0
    PIN CI1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  14.090 1.090 14.170 1.310 ;
        RECT  14.170 1.005 14.310 1.515 ;
        END
    END CI1
    PIN CI0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.750 1.515 ;
        RECT  3.750 1.080 3.960 1.300 ;
        END
    END CI0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.060 3.290 1.280 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.840 0.300 ;
        RECT  6.840 -0.300 6.960 0.520 ;
        RECT  6.960 -0.300 8.235 0.300 ;
        RECT  8.235 -0.300 8.355 0.520 ;
        RECT  8.355 -0.300 9.745 0.300 ;
        RECT  9.745 -0.300 9.865 0.520 ;
        RECT  9.865 -0.300 11.070 0.300 ;
        RECT  11.070 -0.300 11.190 0.520 ;
        RECT  11.190 -0.300 16.915 0.300 ;
        RECT  16.915 -0.300 17.135 0.340 ;
        RECT  17.135 -0.300 17.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 16.915 2.820 ;
        RECT  16.915 2.180 17.135 2.820 ;
        RECT  17.135 2.220 17.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.890 0.730 12.020 1.570 ;
        RECT  12.020 0.730 12.210 0.910 ;
        RECT  2.890 1.050 2.900 2.050 ;
        RECT  2.900 0.760 3.030 2.050 ;
        RECT  3.030 1.470 3.050 2.050 ;
        RECT  3.030 0.760 3.140 0.920 ;
        RECT  3.050 1.930 6.150 2.050 ;
        RECT  6.150 1.930 6.370 2.070 ;
        RECT  6.370 1.930 11.710 2.050 ;
        RECT  11.710 1.930 11.950 2.070 ;
        RECT  11.480 1.090 11.550 1.570 ;
        RECT  11.550 0.720 11.600 1.570 ;
        RECT  11.600 0.720 11.690 1.210 ;
        RECT  11.690 0.990 11.770 1.210 ;
        RECT  10.570 0.720 10.710 1.810 ;
        RECT  10.710 1.670 10.880 1.810 ;
        RECT  7.320 0.720 7.440 1.810 ;
        RECT  7.440 0.720 7.460 1.505 ;
        RECT  7.460 1.345 7.980 1.505 ;
        RECT  5.600 0.710 5.720 1.260 ;
        RECT  5.720 1.120 5.780 1.260 ;
        RECT  5.780 1.120 5.920 1.810 ;
        RECT  5.920 1.690 6.870 1.810 ;
        RECT  6.870 1.180 6.980 1.810 ;
        RECT  6.980 1.060 6.990 1.810 ;
        RECT  6.990 1.060 7.150 1.300 ;
        RECT  6.340 0.720 6.480 1.250 ;
        RECT  6.480 1.130 6.600 1.570 ;
        RECT  6.600 1.430 6.730 1.570 ;
        RECT  6.040 0.730 6.170 1.570 ;
        RECT  6.170 1.430 6.350 1.570 ;
        RECT  3.770 1.690 4.080 1.810 ;
        RECT  3.530 0.710 4.080 0.870 ;
        RECT  4.080 0.710 4.200 1.810 ;
        RECT  4.200 1.050 4.340 1.210 ;
        RECT  5.170 0.710 5.320 1.260 ;
        RECT  4.200 1.690 5.340 1.810 ;
        RECT  5.320 1.120 5.340 1.260 ;
        RECT  5.340 1.120 5.460 1.810 ;
        RECT  5.460 1.120 5.480 1.680 ;
        RECT  5.480 1.520 5.610 1.680 ;
        RECT  2.260 0.470 2.360 0.660 ;
        RECT  2.260 1.590 2.380 1.750 ;
        RECT  2.360 0.470 4.590 0.590 ;
        RECT  4.590 0.420 4.810 0.590 ;
        RECT  4.320 0.760 4.505 0.920 ;
        RECT  4.505 0.760 4.625 1.560 ;
        RECT  0.420 0.480 0.640 0.880 ;
        RECT  0.640 1.895 0.850 2.015 ;
        RECT  0.640 0.760 0.850 0.880 ;
        RECT  0.850 0.760 0.990 2.015 ;
        RECT  0.990 1.090 1.460 1.250 ;
        RECT  0.990 1.895 2.550 2.015 ;
        RECT  2.540 0.710 2.550 0.830 ;
        RECT  2.550 0.710 2.690 2.015 ;
        RECT  2.690 1.470 2.710 2.015 ;
        RECT  2.690 0.710 2.780 0.850 ;
        RECT  1.330 0.780 1.760 0.900 ;
        RECT  1.110 1.570 1.860 1.730 ;
        RECT  1.760 0.480 1.860 0.900 ;
        RECT  1.860 0.480 1.980 1.730 ;
        RECT  12.480 0.710 12.540 0.940 ;
        RECT  12.360 0.710 12.480 1.260 ;
        RECT  12.330 1.120 12.360 1.260 ;
        RECT  12.210 1.120 12.330 1.810 ;
        RECT  12.140 1.590 12.210 1.810 ;
        RECT  11.130 1.690 12.140 1.810 ;
        RECT  11.010 1.080 11.130 1.810 ;
        RECT  13.240 0.740 13.350 0.900 ;
        RECT  13.100 0.740 13.240 1.570 ;
        RECT  13.880 0.740 14.460 0.880 ;
        RECT  13.880 1.670 14.450 1.810 ;
        RECT  13.720 0.740 13.880 1.810 ;
        RECT  12.740 1.690 13.720 1.810 ;
        RECT  12.760 0.710 12.920 1.260 ;
        RECT  12.740 1.120 12.760 1.260 ;
        RECT  12.620 1.120 12.740 1.810 ;
        RECT  12.600 1.120 12.620 1.720 ;
        RECT  14.760 0.710 14.780 0.930 ;
        RECT  14.590 0.710 14.760 2.050 ;
        RECT  13.160 1.930 14.590 2.050 ;
        RECT  15.440 0.420 15.660 0.590 ;
        RECT  15.440 1.590 15.560 1.810 ;
        RECT  15.420 0.470 15.440 1.810 ;
        RECT  15.320 0.470 15.420 1.710 ;
        RECT  11.430 0.470 15.320 0.590 ;
        RECT  11.310 0.470 11.430 0.760 ;
        RECT  10.950 0.640 11.310 0.760 ;
        RECT  10.830 0.470 10.950 0.760 ;
        RECT  10.105 0.470 10.830 0.590 ;
        RECT  9.985 0.470 10.105 0.760 ;
        RECT  9.625 0.640 9.985 0.760 ;
        RECT  9.505 0.470 9.625 0.760 ;
        RECT  8.595 0.470 9.505 0.590 ;
        RECT  8.475 0.470 8.595 0.760 ;
        RECT  8.115 0.640 8.475 0.760 ;
        RECT  7.995 0.470 8.115 0.760 ;
        RECT  7.200 0.470 7.995 0.590 ;
        RECT  7.080 0.470 7.200 0.760 ;
        RECT  6.720 0.640 7.080 0.760 ;
        RECT  6.600 0.470 6.720 0.760 ;
        RECT  5.050 0.470 6.600 0.590 ;
        RECT  5.050 1.430 5.210 1.570 ;
        RECT  4.930 0.470 5.050 1.570 ;
        RECT  4.910 0.740 4.930 1.570 ;
        RECT  15.800 1.495 15.980 1.655 ;
        RECT  15.800 0.720 15.855 0.940 ;
        RECT  15.680 0.720 15.800 1.655 ;
        RECT  16.360 1.080 16.590 1.240 ;
        RECT  16.240 1.080 16.360 2.050 ;
        RECT  15.200 1.930 16.240 2.050 ;
        RECT  15.120 1.890 15.200 2.050 ;
        RECT  15.120 0.710 15.190 0.940 ;
        RECT  15.560 1.030 15.680 1.250 ;
        RECT  4.750 0.740 4.910 0.900 ;
        RECT  12.920 1.930 13.160 2.070 ;
        RECT  12.470 1.560 12.600 1.720 ;
        RECT  12.870 1.430 13.100 1.570 ;
        RECT  10.930 1.080 11.010 1.300 ;
        RECT  11.730 1.430 11.890 1.570 ;
        RECT  2.810 1.050 2.890 1.270 ;
        RECT  11.350 1.430 11.480 1.570 ;
        RECT  9.990 1.345 10.570 1.505 ;
        RECT  7.170 1.670 7.320 1.810 ;
        RECT  14.980 0.710 15.120 2.050 ;
        RECT  5.540 0.710 5.600 0.940 ;
        RECT  6.290 1.030 6.340 1.250 ;
        RECT  5.870 0.730 6.040 0.910 ;
        RECT  3.530 1.670 3.770 1.810 ;
        RECT  2.140 0.470 2.260 1.750 ;
        RECT  4.350 1.400 4.505 1.560 ;
        RECT  0.420 1.595 0.640 2.015 ;
        RECT  1.110 0.480 1.330 0.900 ;
    END
END FCSICOND2

MACRO FICIND1
    CLASS CORE ;
    FOREIGN FICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.650 1.940 7.680 2.100 ;
        RECT  7.680 1.390 7.770 2.100 ;
        RECT  7.680 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.840 2.100 ;
        RECT  7.840 1.940 7.870 2.100 ;
        RECT  7.840 0.780 7.910 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 0.450 6.950 1.550 ;
        RECT  6.950 0.450 7.030 0.900 ;
        RECT  6.950 1.410 7.050 1.550 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.965 2.010 1.185 ;
        RECT  2.010 0.965 2.150 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 7.235 0.300 ;
        RECT  7.235 -0.300 7.455 0.340 ;
        RECT  7.455 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 7.235 2.820 ;
        RECT  7.235 2.180 7.455 2.820 ;
        RECT  7.455 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.170 0.590 4.220 2.050 ;
        RECT  4.220 0.590 4.290 1.750 ;
        RECT  3.740 0.500 3.850 0.920 ;
        RECT  3.850 0.500 3.970 1.810 ;
        RECT  3.970 1.050 4.050 1.270 ;
        RECT  2.400 0.470 2.500 0.630 ;
        RECT  2.400 1.615 2.520 1.775 ;
        RECT  2.500 0.470 3.455 0.590 ;
        RECT  3.455 0.470 3.575 1.270 ;
        RECT  3.575 1.050 3.730 1.270 ;
        RECT  0.560 0.480 0.780 0.880 ;
        RECT  0.780 1.895 0.990 2.015 ;
        RECT  0.780 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.110 2.015 ;
        RECT  1.110 1.080 1.320 1.240 ;
        RECT  1.110 1.895 2.670 2.015 ;
        RECT  2.670 0.710 2.810 2.015 ;
        RECT  2.810 1.470 2.850 2.015 ;
        RECT  2.810 0.710 2.920 0.850 ;
        RECT  1.250 0.480 1.440 0.900 ;
        RECT  1.440 0.480 1.470 1.775 ;
        RECT  1.470 0.570 1.560 1.775 ;
        RECT  1.560 1.635 2.140 1.775 ;
        RECT  1.560 0.570 2.140 0.730 ;
        RECT  4.130 0.590 4.170 0.830 ;
        RECT  4.100 1.530 4.170 2.050 ;
        RECT  3.190 1.930 4.100 2.050 ;
        RECT  3.190 0.760 3.290 0.920 ;
        RECT  3.050 0.760 3.190 2.050 ;
        RECT  3.030 1.050 3.050 2.050 ;
        RECT  6.330 1.050 6.405 1.270 ;
        RECT  6.210 0.710 6.330 1.540 ;
        RECT  5.670 0.710 6.210 0.850 ;
        RECT  6.550 0.470 6.670 1.550 ;
        RECT  6.490 0.470 6.550 0.950 ;
        RECT  6.450 1.410 6.550 1.550 ;
        RECT  5.050 0.470 6.490 0.590 ;
        RECT  4.990 0.470 5.050 0.770 ;
        RECT  4.990 1.410 5.010 1.650 ;
        RECT  6.620 1.910 6.860 2.070 ;
        RECT  4.680 1.910 6.620 2.050 ;
        RECT  4.540 0.590 4.680 2.050 ;
        RECT  4.520 0.590 4.540 1.710 ;
        RECT  7.540 1.060 7.610 1.280 ;
        RECT  7.420 1.060 7.540 1.790 ;
        RECT  5.400 1.670 7.420 1.790 ;
        RECT  5.290 0.710 5.540 0.850 ;
        RECT  5.290 1.430 5.400 1.790 ;
        RECT  5.280 0.710 5.290 1.790 ;
        RECT  4.410 1.550 4.520 1.710 ;
        RECT  4.850 0.470 4.990 1.650 ;
        RECT  5.570 1.400 6.210 1.540 ;
        RECT  2.930 1.050 3.030 1.270 ;
        RECT  5.170 0.710 5.280 1.650 ;
        RECT  3.710 1.410 3.850 1.810 ;
        RECT  2.280 0.470 2.400 1.775 ;
        RECT  0.560 1.595 0.780 2.015 ;
        RECT  1.230 1.615 1.440 1.775 ;
    END
END FICIND1

MACRO FICIND2
    CLASS CORE ;
    FOREIGN FICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 0.750 7.900 1.755 ;
        RECT  7.900 0.450 7.910 1.755 ;
        RECT  7.910 0.450 8.120 0.870 ;
        RECT  7.910 1.595 8.140 1.755 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.130 0.750 7.180 1.550 ;
        RECT  7.180 0.450 7.270 1.550 ;
        RECT  7.270 0.450 7.400 0.870 ;
        RECT  7.270 1.410 7.420 1.550 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END CIN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 0.965 2.010 1.185 ;
        RECT  2.010 0.965 2.150 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 8.290 0.300 ;
        RECT  8.290 -0.300 8.510 0.340 ;
        RECT  8.510 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 8.290 2.820 ;
        RECT  8.290 2.180 8.510 2.820 ;
        RECT  8.510 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.400 0.470 2.500 0.630 ;
        RECT  2.400 1.490 2.520 1.650 ;
        RECT  2.500 0.470 3.455 0.590 ;
        RECT  3.455 0.470 3.575 1.270 ;
        RECT  3.575 1.050 3.730 1.270 ;
        RECT  0.560 0.480 0.780 0.880 ;
        RECT  0.780 1.895 0.990 2.015 ;
        RECT  0.780 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.110 2.015 ;
        RECT  1.110 1.080 1.320 1.240 ;
        RECT  1.110 1.895 2.670 2.015 ;
        RECT  2.670 0.710 2.810 2.015 ;
        RECT  2.810 1.470 2.850 2.015 ;
        RECT  2.810 0.710 2.920 0.850 ;
        RECT  1.250 0.480 1.440 0.900 ;
        RECT  1.440 0.480 1.470 1.775 ;
        RECT  1.470 0.570 1.560 1.775 ;
        RECT  1.560 1.635 2.140 1.775 ;
        RECT  1.560 0.570 2.140 0.730 ;
        RECT  3.970 1.050 4.050 1.270 ;
        RECT  3.930 0.500 3.970 1.530 ;
        RECT  3.850 0.500 3.930 1.810 ;
        RECT  3.740 0.500 3.850 0.920 ;
        RECT  4.220 0.620 4.290 1.750 ;
        RECT  4.170 0.620 4.220 2.050 ;
        RECT  4.130 0.620 4.170 0.860 ;
        RECT  4.100 1.530 4.170 2.050 ;
        RECT  3.190 1.930 4.100 2.050 ;
        RECT  3.190 0.760 3.290 0.920 ;
        RECT  3.050 0.760 3.190 2.050 ;
        RECT  3.030 1.050 3.050 2.050 ;
        RECT  6.330 1.050 6.405 1.270 ;
        RECT  6.210 0.710 6.330 1.540 ;
        RECT  5.670 0.710 6.210 0.850 ;
        RECT  6.650 0.830 6.680 1.550 ;
        RECT  6.560 0.470 6.650 1.550 ;
        RECT  6.490 0.470 6.560 0.950 ;
        RECT  6.450 1.410 6.560 1.550 ;
        RECT  5.050 0.470 6.490 0.590 ;
        RECT  5.010 0.470 5.050 0.770 ;
        RECT  4.910 0.470 5.010 1.650 ;
        RECT  6.620 1.910 6.860 2.070 ;
        RECT  4.680 1.910 6.620 2.050 ;
        RECT  4.540 0.620 4.680 2.050 ;
        RECT  4.520 0.620 4.540 1.710 ;
        RECT  8.260 1.030 8.420 2.050 ;
        RECT  7.330 1.930 8.260 2.050 ;
        RECT  7.210 1.670 7.330 2.050 ;
        RECT  5.400 1.670 7.210 1.790 ;
        RECT  5.290 0.710 5.540 0.850 ;
        RECT  5.290 1.430 5.400 1.790 ;
        RECT  5.280 0.710 5.290 1.790 ;
        RECT  5.170 0.710 5.280 1.650 ;
        RECT  4.410 1.550 4.520 1.710 ;
        RECT  4.850 0.650 4.910 1.650 ;
        RECT  5.570 1.400 6.210 1.540 ;
        RECT  2.930 1.050 3.030 1.270 ;
        RECT  3.710 1.410 3.850 1.810 ;
        RECT  2.280 0.470 2.400 1.650 ;
        RECT  0.560 1.595 0.780 2.015 ;
        RECT  1.230 1.615 1.440 1.775 ;
    END
END FICIND2

MACRO FICOND1
    CLASS CORE ;
    FOREIGN FICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.350 1.940 8.380 2.100 ;
        RECT  8.380 1.390 8.410 2.100 ;
        RECT  8.380 0.420 8.410 0.905 ;
        RECT  8.410 0.420 8.540 2.100 ;
        RECT  8.540 0.785 8.550 1.515 ;
        RECT  8.540 1.940 8.570 2.100 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.540 1.410 7.770 1.550 ;
        RECT  7.560 0.445 7.770 0.870 ;
        RECT  7.770 0.445 7.780 1.550 ;
        RECT  7.780 0.750 7.910 1.550 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.005 6.950 1.235 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.040 2.010 1.260 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.000 0.550 1.515 ;
        RECT  0.550 1.020 0.610 1.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 7.160 0.300 ;
        RECT  7.160 -0.300 7.380 0.340 ;
        RECT  7.380 -0.300 7.935 0.300 ;
        RECT  7.935 -0.300 8.155 0.340 ;
        RECT  8.155 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 7.160 2.820 ;
        RECT  7.160 2.180 7.380 2.820 ;
        RECT  7.380 2.220 7.935 2.820 ;
        RECT  7.935 2.180 8.155 2.820 ;
        RECT  8.155 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.190 0.760 3.290 0.920 ;
        RECT  3.190 1.930 4.100 2.050 ;
        RECT  4.100 1.540 4.170 2.050 ;
        RECT  4.130 0.620 4.170 0.860 ;
        RECT  4.170 0.620 4.220 2.050 ;
        RECT  4.220 0.620 4.290 1.760 ;
        RECT  3.790 0.450 3.850 0.950 ;
        RECT  3.850 0.450 3.970 1.810 ;
        RECT  3.970 1.040 4.050 1.260 ;
        RECT  2.400 0.470 2.500 0.630 ;
        RECT  2.400 1.490 2.520 1.650 ;
        RECT  2.500 0.470 3.550 0.590 ;
        RECT  3.550 0.470 3.670 1.275 ;
        RECT  3.670 1.055 3.730 1.275 ;
        RECT  0.560 0.480 0.780 0.880 ;
        RECT  0.780 1.895 0.985 2.015 ;
        RECT  0.780 0.760 0.985 0.880 ;
        RECT  0.985 0.760 1.105 2.015 ;
        RECT  1.105 1.090 1.270 1.250 ;
        RECT  1.105 1.895 2.690 2.015 ;
        RECT  2.680 0.710 2.690 0.850 ;
        RECT  2.690 0.710 2.830 2.015 ;
        RECT  2.830 1.470 2.850 2.015 ;
        RECT  2.830 0.710 2.920 0.850 ;
        RECT  1.250 0.440 1.405 0.860 ;
        RECT  1.405 0.440 1.470 1.775 ;
        RECT  1.470 0.520 1.525 1.775 ;
        RECT  1.525 1.635 2.140 1.775 ;
        RECT  1.525 0.520 2.140 0.680 ;
        RECT  3.050 0.760 3.190 2.050 ;
        RECT  3.030 1.050 3.050 2.050 ;
        RECT  5.760 0.760 5.950 0.920 ;
        RECT  5.760 1.400 5.850 1.540 ;
        RECT  5.640 0.760 5.760 1.540 ;
        RECT  6.400 0.450 6.620 0.870 ;
        RECT  6.250 1.410 6.610 1.550 ;
        RECT  6.250 0.470 6.400 0.590 ;
        RECT  6.130 0.470 6.250 1.550 ;
        RECT  5.090 0.470 6.130 0.590 ;
        RECT  5.890 1.090 6.130 1.250 ;
        RECT  4.930 0.470 5.090 1.580 ;
        RECT  6.560 1.910 6.800 2.070 ;
        RECT  4.680 1.910 6.560 2.050 ;
        RECT  4.540 0.620 4.680 2.050 ;
        RECT  4.520 0.620 4.540 1.720 ;
        RECT  7.235 1.090 7.550 1.250 ;
        RECT  7.095 0.750 7.235 1.550 ;
        RECT  6.970 0.750 7.095 0.870 ;
        RECT  6.750 1.410 7.095 1.550 ;
        RECT  8.170 1.060 8.290 1.280 ;
        RECT  8.050 1.060 8.170 1.790 ;
        RECT  5.420 1.670 8.050 1.790 ;
        RECT  5.420 0.710 5.520 0.850 ;
        RECT  5.300 0.710 5.420 1.790 ;
        RECT  6.750 0.450 6.970 0.870 ;
        RECT  4.410 1.560 4.520 1.720 ;
        RECT  5.240 1.380 5.300 1.600 ;
        RECT  4.800 1.420 4.930 1.580 ;
        RECT  5.610 1.400 5.640 1.540 ;
        RECT  2.950 1.050 3.030 1.270 ;
        RECT  3.710 1.410 3.850 1.810 ;
        RECT  2.280 0.470 2.400 1.650 ;
        RECT  0.560 1.635 0.780 2.035 ;
        RECT  1.230 1.615 1.405 1.775 ;
    END
END FICOND1

MACRO FICOND2
    CLASS CORE ;
    FOREIGN FICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.940 8.300 2.100 ;
        RECT  8.300 1.390 8.410 2.100 ;
        RECT  8.300 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.460 2.100 ;
        RECT  8.460 1.940 8.490 2.100 ;
        RECT  8.460 0.780 8.550 1.515 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.490 0.445 7.710 0.870 ;
        RECT  7.470 1.410 7.770 1.550 ;
        RECT  7.710 0.750 7.770 0.870 ;
        RECT  7.770 0.750 7.910 1.550 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.005 6.950 1.235 ;
        END
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.840 1.040 2.010 1.260 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.550 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 7.880 0.300 ;
        RECT  7.880 -0.300 8.100 0.340 ;
        RECT  8.100 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 7.880 2.820 ;
        RECT  7.880 2.180 8.100 2.820 ;
        RECT  8.100 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.560 0.480 0.780 0.880 ;
        RECT  0.780 1.895 0.985 2.015 ;
        RECT  0.780 0.760 0.985 0.880 ;
        RECT  0.985 0.760 1.105 2.015 ;
        RECT  1.105 1.080 1.270 1.240 ;
        RECT  1.105 1.895 2.690 2.015 ;
        RECT  2.680 0.710 2.690 0.850 ;
        RECT  2.690 0.710 2.830 2.015 ;
        RECT  2.830 1.470 2.850 2.015 ;
        RECT  2.830 0.710 2.920 0.850 ;
        RECT  1.250 0.440 1.405 0.860 ;
        RECT  1.405 0.440 1.470 1.775 ;
        RECT  1.470 0.520 1.525 1.775 ;
        RECT  1.525 1.635 2.140 1.775 ;
        RECT  1.525 0.520 2.140 0.680 ;
        RECT  3.670 1.055 3.730 1.275 ;
        RECT  3.550 0.470 3.670 1.275 ;
        RECT  2.500 0.470 3.550 0.590 ;
        RECT  2.400 1.490 2.520 1.650 ;
        RECT  2.400 0.470 2.500 0.630 ;
        RECT  3.970 1.040 4.050 1.260 ;
        RECT  3.850 0.450 3.970 1.810 ;
        RECT  3.790 0.450 3.850 0.950 ;
        RECT  4.220 0.620 4.290 1.760 ;
        RECT  4.170 0.620 4.220 2.050 ;
        RECT  4.130 0.620 4.170 0.860 ;
        RECT  4.100 1.540 4.170 2.050 ;
        RECT  3.170 1.930 4.100 2.050 ;
        RECT  3.170 0.760 3.290 0.920 ;
        RECT  3.050 0.760 3.170 2.050 ;
        RECT  3.030 1.050 3.050 2.050 ;
        RECT  5.760 0.760 5.950 0.920 ;
        RECT  5.760 1.400 5.850 1.540 ;
        RECT  5.640 0.760 5.760 1.540 ;
        RECT  6.400 0.450 6.620 0.870 ;
        RECT  6.250 1.410 6.610 1.550 ;
        RECT  6.250 0.470 6.400 0.590 ;
        RECT  6.130 0.470 6.250 1.550 ;
        RECT  5.090 0.470 6.130 0.590 ;
        RECT  5.890 1.080 6.130 1.240 ;
        RECT  4.930 0.470 5.090 1.580 ;
        RECT  6.560 1.910 6.800 2.070 ;
        RECT  4.680 1.910 6.560 2.050 ;
        RECT  4.540 0.620 4.680 2.050 ;
        RECT  4.520 0.620 4.540 1.720 ;
        RECT  7.235 1.080 7.510 1.240 ;
        RECT  7.095 0.750 7.235 1.550 ;
        RECT  6.980 0.750 7.095 0.870 ;
        RECT  6.750 1.410 7.095 1.550 ;
        RECT  8.150 1.050 8.240 1.270 ;
        RECT  8.030 1.050 8.150 1.790 ;
        RECT  5.420 1.670 8.030 1.790 ;
        RECT  5.420 0.710 5.520 0.850 ;
        RECT  5.300 0.710 5.420 1.790 ;
        RECT  5.240 1.380 5.300 1.600 ;
        RECT  6.750 0.450 6.980 0.870 ;
        RECT  4.410 1.560 4.520 1.720 ;
        RECT  4.800 1.420 4.930 1.580 ;
        RECT  5.610 1.400 5.640 1.540 ;
        RECT  2.950 1.050 3.030 1.270 ;
        RECT  3.710 1.410 3.850 1.810 ;
        RECT  2.280 0.470 2.400 1.650 ;
        RECT  0.560 1.595 0.780 2.015 ;
        RECT  1.230 1.615 1.405 1.775 ;
    END
END FICOND2

MACRO FIICOND1
    CLASS CORE ;
    FOREIGN FIICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.010 1.940 8.040 2.100 ;
        RECT  8.040 1.390 8.090 2.100 ;
        RECT  8.040 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.200 2.100 ;
        RECT  8.200 1.940 8.230 2.100 ;
        RECT  8.200 0.780 8.230 1.515 ;
        END
    END S
    PIN CON1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.710 1.370 0.870 ;
        RECT  1.370 0.710 1.510 1.755 ;
        RECT  1.510 1.595 1.760 1.755 ;
        END
    END CON1
    PIN CON0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.780 0.200 1.510 ;
        RECT  0.200 0.420 0.230 1.510 ;
        RECT  0.230 0.420 0.360 0.900 ;
        RECT  0.560 1.940 0.590 2.100 ;
        RECT  0.230 1.390 0.590 1.510 ;
        RECT  0.590 1.390 0.750 2.100 ;
        RECT  0.750 1.940 0.780 2.100 ;
        END
    END CON0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.130 1.005 7.270 1.515 ;
        RECT  7.270 1.080 7.395 1.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.030 1.210 2.050 ;
        RECT  1.210 1.930 4.450 2.050 ;
        RECT  4.450 1.930 4.690 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.730 1.270 ;
        RECT  0.730 0.470 0.870 1.270 ;
        RECT  0.870 0.470 1.750 0.590 ;
        RECT  1.750 0.470 1.910 1.290 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.820 0.300 ;
        RECT  0.820 -0.300 1.040 0.340 ;
        RECT  1.040 -0.300 1.645 0.300 ;
        RECT  1.645 -0.300 1.865 0.340 ;
        RECT  1.865 -0.300 7.570 0.300 ;
        RECT  7.570 -0.300 7.790 0.340 ;
        RECT  7.790 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 7.570 2.820 ;
        RECT  7.570 2.180 7.790 2.820 ;
        RECT  7.790 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.530 1.940 5.560 2.100 ;
        RECT  5.530 0.780 5.560 1.515 ;
        RECT  5.560 1.050 5.620 1.270 ;
        RECT  4.010 1.670 4.110 1.810 ;
        RECT  4.010 0.710 4.110 0.870 ;
        RECT  4.110 1.690 5.000 1.810 ;
        RECT  5.000 1.050 5.120 1.810 ;
        RECT  5.120 1.050 5.290 1.270 ;
        RECT  4.620 0.470 4.740 1.570 ;
        RECT  4.740 0.470 4.840 0.890 ;
        RECT  4.740 1.410 4.860 1.570 ;
        RECT  2.275 1.595 2.410 1.755 ;
        RECT  2.275 1.080 3.200 1.240 ;
        RECT  2.275 0.470 4.230 0.590 ;
        RECT  4.230 0.470 4.350 1.570 ;
        RECT  4.350 0.470 4.470 0.690 ;
        RECT  4.350 1.410 4.500 1.570 ;
        RECT  2.840 0.720 3.530 0.880 ;
        RECT  3.530 0.720 3.690 1.810 ;
        RECT  3.690 1.650 3.730 1.810 ;
        RECT  5.440 0.420 5.530 2.100 ;
        RECT  5.370 0.420 5.440 0.900 ;
        RECT  5.370 1.390 5.440 2.100 ;
        RECT  5.340 1.940 5.370 2.100 ;
        RECT  6.550 0.750 6.710 0.910 ;
        RECT  6.550 1.590 6.710 1.750 ;
        RECT  6.975 0.710 7.400 0.870 ;
        RECT  7.160 1.640 7.380 2.050 ;
        RECT  6.975 1.930 7.160 2.050 ;
        RECT  6.855 0.710 6.975 2.050 ;
        RECT  6.850 0.710 6.855 1.270 ;
        RECT  5.920 1.930 6.855 2.050 ;
        RECT  6.710 1.045 6.850 1.270 ;
        RECT  5.800 0.730 5.920 2.050 ;
        RECT  5.680 0.730 5.800 0.890 ;
        RECT  7.790 1.050 7.940 1.270 ;
        RECT  7.670 0.470 7.790 1.270 ;
        RECT  6.310 0.470 7.670 0.590 ;
        RECT  6.200 0.470 6.310 0.870 ;
        RECT  6.200 1.650 6.300 1.810 ;
        RECT  6.190 0.470 6.200 1.810 ;
        RECT  5.680 1.735 5.800 1.895 ;
        RECT  6.430 0.750 6.550 1.750 ;
        RECT  3.890 0.710 4.010 1.810 ;
        RECT  4.475 1.070 4.620 1.290 ;
        RECT  2.115 0.470 2.275 1.755 ;
        RECT  6.080 0.710 6.190 1.810 ;
        RECT  2.840 1.650 3.530 1.810 ;
    END
END FIICOND1

MACRO FIICOND2
    CLASS CORE ;
    FOREIGN FIICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.175 1.940 9.205 2.100 ;
        RECT  9.205 1.390 9.365 2.100 ;
        RECT  9.200 0.420 9.365 0.900 ;
        RECT  9.365 1.390 9.370 1.515 ;
        RECT  9.365 0.780 9.370 0.900 ;
        RECT  9.365 1.940 9.395 2.100 ;
        RECT  9.370 0.780 9.510 1.515 ;
        END
    END S
    PIN CON1
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 0.710 2.150 1.755 ;
        RECT  2.150 0.710 2.180 0.930 ;
        RECT  2.150 1.595 2.590 1.755 ;
        RECT  2.590 0.710 2.710 1.755 ;
        RECT  2.710 0.710 2.920 0.870 ;
        END
    END CON1
    PIN CON0
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.430 0.730 1.670 ;
        RECT  0.730 0.800 0.750 1.670 ;
        RECT  0.750 0.800 0.870 1.550 ;
        RECT  0.870 0.800 0.970 0.920 ;
        RECT  0.970 0.420 1.130 0.920 ;
        RECT  0.870 1.430 1.350 1.550 ;
        RECT  1.350 1.430 1.510 1.670 ;
        END
    END CON0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.410 1.005 8.550 1.515 ;
        RECT  8.550 1.080 8.680 1.240 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.080 0.230 2.050 ;
        RECT  0.230 1.080 0.610 1.240 ;
        RECT  0.230 1.930 1.680 2.050 ;
        RECT  1.680 1.030 1.840 2.050 ;
        RECT  1.840 1.930 2.850 2.050 ;
        RECT  2.850 1.030 3.005 2.050 ;
        RECT  3.005 1.930 5.735 2.050 ;
        RECT  5.735 1.930 5.975 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.050 1.370 1.270 ;
        RECT  1.370 0.470 1.520 1.270 ;
        RECT  1.520 0.470 2.330 0.590 ;
        RECT  2.330 0.470 2.470 1.290 ;
        RECT  2.470 0.470 3.150 0.590 ;
        RECT  3.150 0.470 3.270 1.240 ;
        RECT  3.270 1.080 3.420 1.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.235 0.300 ;
        RECT  0.235 -0.300 0.455 0.340 ;
        RECT  0.455 -0.300 9.570 0.300 ;
        RECT  9.570 -0.300 9.790 0.340 ;
        RECT  9.790 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 9.570 2.820 ;
        RECT  9.570 2.180 9.790 2.820 ;
        RECT  9.790 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.295 1.670 5.395 1.810 ;
        RECT  5.295 0.710 5.395 0.870 ;
        RECT  5.395 1.690 6.285 1.810 ;
        RECT  6.285 1.050 6.405 1.810 ;
        RECT  6.405 1.050 6.575 1.270 ;
        RECT  5.905 0.470 6.025 1.570 ;
        RECT  6.025 0.470 6.125 0.890 ;
        RECT  6.025 1.410 6.145 1.570 ;
        RECT  3.400 0.470 3.555 0.950 ;
        RECT  3.555 0.470 3.675 1.755 ;
        RECT  3.675 1.080 4.485 1.240 ;
        RECT  3.675 0.470 5.515 0.590 ;
        RECT  5.515 0.470 5.635 1.570 ;
        RECT  5.635 0.470 5.755 0.690 ;
        RECT  5.635 1.410 5.785 1.570 ;
        RECT  4.125 0.720 4.815 0.880 ;
        RECT  4.815 0.720 4.975 1.810 ;
        RECT  4.975 1.650 5.015 1.810 ;
        RECT  6.845 1.050 6.905 1.270 ;
        RECT  6.815 0.780 6.845 1.510 ;
        RECT  6.815 1.940 6.845 2.100 ;
        RECT  6.725 0.420 6.815 2.100 ;
        RECT  6.650 0.420 6.725 0.900 ;
        RECT  6.655 1.390 6.725 2.100 ;
        RECT  7.835 0.750 7.995 0.910 ;
        RECT  7.835 1.590 7.995 1.750 ;
        RECT  8.260 0.710 8.685 0.870 ;
        RECT  8.445 1.640 8.665 2.050 ;
        RECT  8.260 1.930 8.445 2.050 ;
        RECT  8.140 0.710 8.260 2.050 ;
        RECT  8.135 0.710 8.140 1.270 ;
        RECT  7.205 1.930 8.140 2.050 ;
        RECT  7.995 1.045 8.135 1.270 ;
        RECT  7.085 0.730 7.205 2.050 ;
        RECT  6.965 0.730 7.085 0.890 ;
        RECT  9.000 1.050 9.185 1.270 ;
        RECT  8.880 0.470 9.000 1.270 ;
        RECT  7.595 0.470 8.880 0.590 ;
        RECT  7.485 0.470 7.595 0.870 ;
        RECT  7.485 1.650 7.585 1.810 ;
        RECT  7.475 0.470 7.485 1.810 ;
        RECT  6.965 1.735 7.085 1.895 ;
        RECT  7.715 0.750 7.835 1.750 ;
        RECT  7.365 0.710 7.475 1.810 ;
        RECT  6.625 1.940 6.655 2.100 ;
        RECT  5.175 0.710 5.295 1.810 ;
        RECT  5.760 1.070 5.905 1.290 ;
        RECT  3.435 1.595 3.555 1.755 ;
        RECT  4.125 1.650 4.815 1.810 ;
    END
END FIICOND2

MACRO FILL1
    CLASS CORE ;
    FOREIGN FILL1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.320 2.820 ;
        END
    END VDD
END FILL1

MACRO FILL16
    CLASS CORE ;
    FOREIGN FILL16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.140 0.320 ;
        RECT  1.140 -0.300 2.160 0.300 ;
        RECT  2.160 -0.300 2.420 0.320 ;
        RECT  2.420 -0.300 3.440 0.300 ;
        RECT  3.440 -0.300 3.700 0.320 ;
        RECT  3.700 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.980 0.320 ;
        RECT  4.980 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.120 2.820 ;
        END
    END VDD
END FILL16

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
END FILL2

MACRO FILL32
    CLASS CORE ;
    FOREIGN FILL32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.140 0.320 ;
        RECT  1.140 -0.300 2.160 0.300 ;
        RECT  2.160 -0.300 2.420 0.320 ;
        RECT  2.420 -0.300 3.440 0.300 ;
        RECT  3.440 -0.300 3.700 0.320 ;
        RECT  3.700 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.980 0.320 ;
        RECT  4.980 -0.300 6.000 0.300 ;
        RECT  6.000 -0.300 6.260 0.320 ;
        RECT  6.260 -0.300 7.280 0.300 ;
        RECT  7.280 -0.300 7.540 0.320 ;
        RECT  7.540 -0.300 8.560 0.300 ;
        RECT  8.560 -0.300 8.820 0.320 ;
        RECT  8.820 -0.300 9.840 0.300 ;
        RECT  9.840 -0.300 10.100 0.320 ;
        RECT  10.100 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 10.240 2.820 ;
        END
    END VDD
END FILL32

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.140 0.320 ;
        RECT  1.140 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.280 2.820 ;
        END
    END VDD
END FILL4

MACRO FILL64
    CLASS CORE ;
    FOREIGN FILL64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.140 0.320 ;
        RECT  1.140 -0.300 2.160 0.300 ;
        RECT  2.160 -0.300 2.420 0.320 ;
        RECT  2.420 -0.300 3.440 0.300 ;
        RECT  3.440 -0.300 3.700 0.320 ;
        RECT  3.700 -0.300 4.720 0.300 ;
        RECT  4.720 -0.300 4.980 0.320 ;
        RECT  4.980 -0.300 6.000 0.300 ;
        RECT  6.000 -0.300 6.260 0.320 ;
        RECT  6.260 -0.300 7.280 0.300 ;
        RECT  7.280 -0.300 7.540 0.320 ;
        RECT  7.540 -0.300 8.560 0.300 ;
        RECT  8.560 -0.300 8.820 0.320 ;
        RECT  8.820 -0.300 9.840 0.300 ;
        RECT  9.840 -0.300 10.100 0.320 ;
        RECT  10.100 -0.300 11.120 0.300 ;
        RECT  11.120 -0.300 11.380 0.320 ;
        RECT  11.380 -0.300 12.400 0.300 ;
        RECT  12.400 -0.300 12.660 0.320 ;
        RECT  12.660 -0.300 13.680 0.300 ;
        RECT  13.680 -0.300 13.940 0.320 ;
        RECT  13.940 -0.300 14.960 0.300 ;
        RECT  14.960 -0.300 15.220 0.320 ;
        RECT  15.220 -0.300 16.240 0.300 ;
        RECT  16.240 -0.300 16.500 0.320 ;
        RECT  16.500 -0.300 17.520 0.300 ;
        RECT  17.520 -0.300 17.780 0.320 ;
        RECT  17.780 -0.300 18.800 0.300 ;
        RECT  18.800 -0.300 19.060 0.320 ;
        RECT  19.060 -0.300 20.080 0.300 ;
        RECT  20.080 -0.300 20.340 0.320 ;
        RECT  20.340 -0.300 20.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 20.480 2.820 ;
        END
    END VDD
END FILL64

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.880 0.300 ;
        RECT  0.880 -0.300 1.140 0.320 ;
        RECT  1.140 -0.300 2.160 0.300 ;
        RECT  2.160 -0.300 2.420 0.320 ;
        RECT  2.420 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
END FILL8

MACRO HA1D1
    CLASS CORE ;
    FOREIGN HA1D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.960 4.230 2.100 ;
        RECT  4.230 1.390 4.250 2.100 ;
        RECT  4.230 0.420 4.250 0.955 ;
        RECT  4.250 0.420 4.390 2.100 ;
        RECT  4.390 1.960 4.420 2.100 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.060 1.960 0.080 2.100 ;
        RECT  0.080 0.420 0.200 2.100 ;
        RECT  0.200 1.390 0.250 2.100 ;
        RECT  0.200 0.420 0.250 0.955 ;
        RECT  0.250 1.960 0.280 2.100 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.360 1.160 1.515 ;
        RECT  1.160 1.360 1.280 2.050 ;
        RECT  1.280 1.930 3.410 2.050 ;
        RECT  3.410 1.930 3.650 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.210 2.820 ;
        RECT  1.210 2.180 1.430 2.820 ;
        RECT  1.430 2.220 1.990 2.820 ;
        RECT  1.990 2.180 2.210 2.820 ;
        RECT  2.210 2.220 3.800 2.820 ;
        RECT  3.800 2.180 4.020 2.820 ;
        RECT  4.020 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.990 1.030 4.110 1.810 ;
        RECT  4.110 1.030 4.130 1.270 ;
        RECT  3.490 0.590 3.610 1.570 ;
        RECT  3.610 1.410 3.730 1.570 ;
        RECT  3.610 0.590 3.730 0.750 ;
        RECT  1.700 0.470 1.920 0.885 ;
        RECT  1.820 1.410 2.090 1.530 ;
        RECT  1.920 0.470 2.090 0.590 ;
        RECT  2.090 0.470 2.230 1.530 ;
        RECT  2.230 1.050 2.370 1.270 ;
        RECT  2.230 0.470 3.140 0.590 ;
        RECT  3.140 0.470 3.260 1.570 ;
        RECT  3.260 1.410 3.370 1.570 ;
        RECT  3.260 0.650 3.370 0.810 ;
        RECT  2.370 0.710 2.490 0.850 ;
        RECT  2.490 0.710 2.610 1.810 ;
        RECT  0.380 0.750 0.500 1.760 ;
        RECT  0.500 1.640 0.820 1.760 ;
        RECT  0.820 1.640 1.040 2.060 ;
        RECT  0.500 0.750 1.060 0.870 ;
        RECT  1.060 0.450 1.280 0.870 ;
        RECT  2.980 1.690 3.990 1.810 ;
        RECT  2.850 0.710 3.010 0.850 ;
        RECT  2.850 1.640 2.980 1.810 ;
        RECT  2.730 0.710 2.850 1.810 ;
        RECT  3.380 1.040 3.490 1.200 ;
        RECT  1.600 1.410 1.820 1.810 ;
        RECT  2.380 1.410 2.490 1.810 ;
        RECT  0.320 1.055 0.380 1.275 ;
    END
END HA1D1

MACRO HA1D2
    CLASS CORE ;
    FOREIGN HA1D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.960 4.510 2.100 ;
        RECT  4.510 1.390 4.570 2.100 ;
        RECT  4.510 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.670 2.100 ;
        RECT  4.670 1.960 4.700 2.100 ;
        RECT  4.670 0.780 4.710 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.470 0.230 2.040 ;
        RECT  0.230 1.880 0.660 2.040 ;
        RECT  0.230 0.470 0.660 0.630 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.360 1.460 1.515 ;
        RECT  1.460 1.360 1.580 2.050 ;
        RECT  1.580 1.930 3.710 2.050 ;
        RECT  3.710 1.930 3.950 2.090 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 2.290 2.820 ;
        RECT  2.290 2.180 2.510 2.820 ;
        RECT  2.510 2.220 4.080 2.820 ;
        RECT  4.080 2.180 4.300 2.820 ;
        RECT  4.300 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.800 0.750 1.360 0.870 ;
        RECT  1.360 0.450 1.580 0.870 ;
        RECT  1.120 1.640 1.340 2.060 ;
        RECT  0.800 1.640 1.120 1.760 ;
        RECT  0.680 0.750 0.800 1.760 ;
        RECT  2.790 0.710 2.910 1.810 ;
        RECT  2.670 0.710 2.790 0.850 ;
        RECT  3.560 0.650 3.670 0.810 ;
        RECT  3.560 1.410 3.670 1.570 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  2.530 0.470 3.440 0.590 ;
        RECT  2.530 1.050 2.670 1.270 ;
        RECT  2.390 0.470 2.530 1.530 ;
        RECT  2.220 0.470 2.390 0.590 ;
        RECT  2.120 1.410 2.390 1.530 ;
        RECT  2.000 0.470 2.220 0.885 ;
        RECT  3.910 0.590 4.030 0.750 ;
        RECT  3.910 1.410 4.030 1.570 ;
        RECT  3.790 0.590 3.910 1.570 ;
        RECT  4.390 1.030 4.450 1.270 ;
        RECT  4.270 1.030 4.390 1.810 ;
        RECT  3.280 1.690 4.270 1.810 ;
        RECT  3.150 0.710 3.310 0.850 ;
        RECT  3.150 1.640 3.280 1.810 ;
        RECT  3.680 1.040 3.790 1.200 ;
        RECT  1.900 1.410 2.120 1.810 ;
        RECT  2.680 1.410 2.790 1.810 ;
        RECT  0.400 1.080 0.680 1.240 ;
        RECT  3.030 0.710 3.150 1.810 ;
    END
END HA1D2

MACRO HA1D4
    CLASS CORE ;
    FOREIGN HA1D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.990 1.650 7.310 2.030 ;
        RECT  6.990 0.490 7.310 0.870 ;
        RECT  7.310 0.490 7.730 2.030 ;
        RECT  7.730 1.650 7.910 2.030 ;
        RECT  7.730 0.490 7.910 0.870 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.650 0.590 2.030 ;
        RECT  0.420 0.490 0.590 0.870 ;
        RECT  0.590 0.490 1.010 2.030 ;
        RECT  1.010 1.650 1.330 2.030 ;
        RECT  1.010 0.490 1.330 0.870 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.080 2.010 1.240 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.395 2.780 1.515 ;
        RECT  2.780 1.050 2.870 1.515 ;
        RECT  2.870 1.050 2.940 2.050 ;
        RECT  2.940 1.360 2.990 2.050 ;
        RECT  2.990 1.930 6.150 2.050 ;
        RECT  6.150 1.930 6.390 2.070 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.080 2.540 1.240 ;
        RECT  2.540 0.810 2.660 1.240 ;
        RECT  2.660 0.810 3.290 0.930 ;
        RECT  3.290 0.810 3.410 1.235 ;
        RECT  3.410 1.005 3.750 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.530 0.300 ;
        RECT  1.530 -0.300 1.750 0.340 ;
        RECT  1.750 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.060 0.340 ;
        RECT  3.060 -0.300 3.640 0.300 ;
        RECT  3.640 -0.300 3.860 0.340 ;
        RECT  3.860 -0.300 4.800 0.300 ;
        RECT  4.800 -0.300 5.020 0.340 ;
        RECT  5.020 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.640 2.820 ;
        RECT  3.640 2.180 3.860 2.820 ;
        RECT  3.860 2.220 4.790 2.820 ;
        RECT  4.790 2.180 5.010 2.820 ;
        RECT  5.010 2.220 6.590 2.820 ;
        RECT  6.590 2.180 6.810 2.820 ;
        RECT  6.810 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.530 1.635 2.750 2.055 ;
        RECT  2.060 1.635 2.530 1.755 ;
        RECT  2.190 0.430 2.410 0.850 ;
        RECT  1.570 0.730 2.190 0.850 ;
        RECT  1.840 1.635 2.060 2.055 ;
        RECT  1.570 1.635 1.840 1.755 ;
        RECT  1.450 0.730 1.570 1.755 ;
        RECT  5.300 0.710 5.420 1.810 ;
        RECT  4.380 0.710 5.300 0.850 ;
        RECT  5.190 1.410 5.300 1.810 ;
        RECT  4.620 1.690 5.190 1.810 ;
        RECT  6.040 0.660 6.200 0.820 ;
        RECT  6.040 1.410 6.180 1.570 ;
        RECT  5.920 0.470 6.040 1.570 ;
        RECT  4.260 0.470 5.920 0.590 ;
        RECT  4.260 1.080 4.880 1.240 ;
        RECT  4.120 0.470 4.260 1.810 ;
        RECT  3.220 0.470 4.120 0.630 ;
        RECT  4.040 1.410 4.120 1.810 ;
        RECT  3.460 1.410 4.040 1.550 ;
        RECT  6.420 1.410 6.540 1.570 ;
        RECT  6.420 0.660 6.490 1.240 ;
        RECT  6.330 0.660 6.420 1.570 ;
        RECT  6.300 1.080 6.330 1.570 ;
        RECT  6.830 1.080 7.095 1.240 ;
        RECT  6.710 1.080 6.830 1.810 ;
        RECT  5.790 1.690 6.710 1.810 ;
        RECT  5.690 0.710 5.800 0.850 ;
        RECT  5.690 1.640 5.790 1.810 ;
        RECT  6.160 1.080 6.300 1.240 ;
        RECT  3.240 1.410 3.460 1.810 ;
        RECT  5.570 0.710 5.690 1.810 ;
        RECT  4.390 1.410 4.620 1.810 ;
        RECT  1.225 1.080 1.450 1.240 ;
        LAYER M1 ;
        RECT  1.225 0.490 1.330 0.870 ;
        RECT  1.225 1.650 1.330 2.030 ;
        RECT  6.990 0.490 7.095 0.870 ;
        RECT  6.990 1.650 7.095 2.030 ;
    END
END HA1D4

MACRO HCOSCIND1
    CLASS CORE ;
    FOREIGN HCOSCIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.040 1.940 8.070 2.100 ;
        RECT  8.070 1.390 8.090 2.100 ;
        RECT  8.070 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.230 2.100 ;
        RECT  8.230 1.940 8.260 2.100 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.330 1.515 ;
        END
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.060 1.940 0.090 2.100 ;
        RECT  0.090 0.420 0.210 2.100 ;
        RECT  0.210 1.390 0.250 2.100 ;
        RECT  0.210 0.420 0.250 0.905 ;
        RECT  0.250 1.940 0.280 2.100 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.140 1.005 5.210 1.230 ;
        RECT  5.210 1.005 5.350 1.515 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.530 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.165 2.820 ;
        RECT  1.165 2.180 1.385 2.820 ;
        RECT  1.385 2.220 2.010 2.820 ;
        RECT  2.010 2.030 2.230 2.820 ;
        RECT  2.230 2.220 2.850 2.820 ;
        RECT  2.850 2.030 3.070 2.820 ;
        RECT  3.070 2.220 5.210 2.820 ;
        RECT  5.210 1.980 5.370 2.820 ;
        RECT  5.370 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.330 1.930 4.190 2.050 ;
        RECT  4.190 1.930 4.410 2.070 ;
        RECT  4.410 1.930 4.900 2.050 ;
        RECT  4.900 0.710 5.020 2.050 ;
        RECT  5.020 1.470 5.090 1.690 ;
        RECT  5.020 0.710 5.160 0.870 ;
        RECT  4.170 0.660 4.230 1.140 ;
        RECT  4.230 0.660 4.350 1.560 ;
        RECT  4.350 1.420 4.470 1.560 ;
        RECT  1.640 0.450 1.740 0.870 ;
        RECT  1.740 0.450 1.860 1.570 ;
        RECT  1.860 1.080 2.730 1.240 ;
        RECT  1.860 0.470 3.740 0.590 ;
        RECT  3.740 0.470 3.860 1.380 ;
        RECT  3.860 1.260 3.920 1.380 ;
        RECT  3.860 0.630 4.020 0.790 ;
        RECT  3.920 1.260 4.080 1.570 ;
        RECT  2.340 0.720 3.030 0.880 ;
        RECT  3.030 0.720 3.190 1.560 ;
        RECT  3.190 1.400 3.350 1.560 ;
        RECT  0.400 0.470 0.520 1.760 ;
        RECT  0.520 1.620 0.750 1.760 ;
        RECT  0.750 1.620 0.970 2.040 ;
        RECT  0.520 0.470 1.000 0.590 ;
        RECT  1.000 0.450 1.220 0.870 ;
        RECT  3.210 1.760 3.330 2.050 ;
        RECT  1.210 1.760 3.210 1.880 ;
        RECT  1.090 1.370 1.210 1.880 ;
        RECT  0.850 1.370 1.090 1.490 ;
        RECT  6.230 0.710 6.470 0.880 ;
        RECT  5.800 1.700 6.470 1.860 ;
        RECT  5.800 0.760 6.230 0.880 ;
        RECT  5.700 0.760 5.800 0.920 ;
        RECT  5.700 1.440 5.800 1.860 ;
        RECT  7.080 0.700 7.230 0.860 ;
        RECT  7.080 1.390 7.180 1.810 ;
        RECT  7.020 0.470 7.080 1.810 ;
        RECT  6.960 0.470 7.020 1.510 ;
        RECT  4.730 0.470 6.960 0.590 ;
        RECT  4.610 0.470 4.730 1.810 ;
        RECT  3.720 1.690 4.610 1.810 ;
        RECT  3.620 1.640 3.720 1.810 ;
        RECT  3.500 0.710 3.620 1.810 ;
        RECT  7.360 0.570 7.520 1.720 ;
        RECT  7.860 1.050 7.970 1.270 ;
        RECT  7.720 1.050 7.860 2.050 ;
        RECT  6.800 1.930 7.720 2.050 ;
        RECT  6.720 0.710 6.830 0.860 ;
        RECT  6.720 1.660 6.800 2.050 ;
        RECT  7.200 1.090 7.360 1.250 ;
        RECT  3.380 0.710 3.500 0.850 ;
        RECT  5.580 0.760 5.700 1.860 ;
        RECT  0.690 1.180 0.850 1.490 ;
        RECT  6.600 0.710 6.720 2.050 ;
        RECT  4.000 0.980 4.170 1.140 ;
        RECT  1.570 1.410 1.740 1.570 ;
        RECT  2.390 1.400 3.030 1.560 ;
        RECT  0.330 1.050 0.400 1.270 ;
    END
END HCOSCIND1

MACRO HCOSCIND2
    CLASS CORE ;
    FOREIGN HCOSCIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.640 1.940 8.670 2.100 ;
        RECT  8.670 1.390 8.730 2.100 ;
        RECT  8.670 0.420 8.730 0.900 ;
        RECT  8.730 0.420 8.830 2.100 ;
        RECT  8.830 1.940 8.860 2.100 ;
        RECT  8.830 0.780 8.870 1.515 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 1.005 6.630 1.515 ;
        RECT  6.630 1.180 6.830 1.400 ;
        END
    END CS
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.785 0.230 1.515 ;
        RECT  0.560 1.940 0.590 2.100 ;
        RECT  0.230 1.390 0.590 1.515 ;
        RECT  0.230 0.785 0.590 0.905 ;
        RECT  0.590 1.390 0.750 2.100 ;
        RECT  0.590 0.420 0.750 0.905 ;
        RECT  0.750 1.940 0.780 2.100 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.640 1.005 5.850 1.230 ;
        RECT  5.850 1.005 5.990 1.515 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 2.150 1.235 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.145 0.300 ;
        RECT  0.145 -0.300 0.365 0.340 ;
        RECT  0.365 -0.300 5.030 0.300 ;
        RECT  5.030 -0.300 5.250 0.340 ;
        RECT  5.250 -0.300 8.230 0.300 ;
        RECT  8.230 -0.300 8.450 0.340 ;
        RECT  8.450 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 1.665 2.820 ;
        RECT  1.665 2.180 1.885 2.820 ;
        RECT  1.885 2.220 2.510 2.820 ;
        RECT  2.510 2.030 2.730 2.820 ;
        RECT  2.730 2.220 3.350 2.820 ;
        RECT  3.350 2.030 3.570 2.820 ;
        RECT  3.570 2.220 5.680 2.820 ;
        RECT  5.680 2.030 5.900 2.820 ;
        RECT  5.900 2.220 6.480 2.820 ;
        RECT  6.480 2.180 6.700 2.820 ;
        RECT  6.700 2.220 8.230 2.820 ;
        RECT  8.230 2.180 8.450 2.820 ;
        RECT  8.450 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.690 1.400 3.850 1.560 ;
        RECT  0.950 0.470 1.070 1.760 ;
        RECT  1.070 1.620 1.250 1.760 ;
        RECT  1.250 1.620 1.470 2.040 ;
        RECT  1.070 0.470 1.500 0.590 ;
        RECT  1.500 0.450 1.720 0.870 ;
        RECT  3.530 0.720 3.690 1.560 ;
        RECT  2.840 0.720 3.530 0.880 ;
        RECT  4.420 1.260 4.580 1.570 ;
        RECT  4.360 0.630 4.520 0.790 ;
        RECT  4.360 1.260 4.420 1.380 ;
        RECT  4.240 0.470 4.360 1.380 ;
        RECT  2.390 0.470 4.240 0.590 ;
        RECT  2.390 1.080 3.230 1.240 ;
        RECT  2.270 0.450 2.390 1.570 ;
        RECT  2.140 0.450 2.270 0.870 ;
        RECT  4.830 1.420 4.970 1.560 ;
        RECT  4.710 0.660 4.830 1.560 ;
        RECT  4.670 0.660 4.710 1.140 ;
        RECT  5.520 0.710 5.660 0.870 ;
        RECT  5.520 1.480 5.590 1.700 ;
        RECT  5.400 0.710 5.520 2.050 ;
        RECT  4.910 1.930 5.400 2.050 ;
        RECT  4.690 1.930 4.910 2.070 ;
        RECT  3.830 1.930 4.690 2.050 ;
        RECT  3.710 1.760 3.830 2.050 ;
        RECT  1.710 1.760 3.710 1.880 ;
        RECT  1.590 1.370 1.710 1.880 ;
        RECT  1.350 1.370 1.590 1.490 ;
        RECT  6.270 0.710 6.970 0.880 ;
        RECT  6.270 1.700 6.970 1.860 ;
        RECT  7.580 0.700 7.730 0.860 ;
        RECT  7.580 1.390 7.680 1.810 ;
        RECT  7.520 0.470 7.580 1.810 ;
        RECT  7.460 0.470 7.520 1.510 ;
        RECT  5.230 0.470 7.460 0.590 ;
        RECT  5.110 0.470 5.230 1.810 ;
        RECT  4.220 1.690 5.110 1.810 ;
        RECT  4.120 1.640 4.220 1.810 ;
        RECT  4.000 0.710 4.120 1.810 ;
        RECT  7.860 0.620 8.020 1.720 ;
        RECT  8.460 1.050 8.570 1.270 ;
        RECT  8.320 1.050 8.460 2.050 ;
        RECT  7.300 1.930 8.320 2.050 ;
        RECT  7.220 0.710 7.330 0.860 ;
        RECT  7.220 1.660 7.300 2.050 ;
        RECT  7.100 0.710 7.220 2.050 ;
        RECT  7.700 1.090 7.860 1.250 ;
        RECT  3.880 0.710 4.000 0.850 ;
        RECT  6.110 0.710 6.270 1.860 ;
        RECT  1.190 1.180 1.350 1.490 ;
        RECT  4.500 0.980 4.670 1.140 ;
        RECT  2.070 1.410 2.270 1.570 ;
        RECT  2.890 1.400 3.530 1.560 ;
        RECT  0.690 1.080 0.950 1.240 ;
    END
END HCOSCIND2

MACRO HCOSCOND1
    CLASS CORE ;
    FOREIGN HCOSCOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.080 1.940 7.110 2.100 ;
        RECT  7.110 1.390 7.130 2.100 ;
        RECT  7.110 0.420 7.130 0.900 ;
        RECT  7.130 0.420 7.270 2.100 ;
        RECT  7.270 1.940 7.300 2.100 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.370 1.515 ;
        END
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.430 1.530 ;
        RECT  0.430 0.725 0.550 1.810 ;
        RECT  0.550 1.410 0.650 1.810 ;
        RECT  0.550 0.725 0.680 0.870 ;
        RECT  0.680 0.450 0.900 0.870 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 2.050 ;
        RECT  0.250 1.930 1.350 2.050 ;
        RECT  1.350 1.760 1.470 2.050 ;
        RECT  1.470 1.760 2.860 1.880 ;
        RECT  2.860 1.760 2.980 2.050 ;
        RECT  2.980 1.930 3.870 2.050 ;
        RECT  3.870 1.930 4.090 2.070 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 1.190 1.240 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.230 0.300 ;
        RECT  4.230 -0.300 4.450 0.340 ;
        RECT  4.450 -0.300 5.020 0.300 ;
        RECT  5.020 -0.300 5.240 0.340 ;
        RECT  5.240 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.830 2.820 ;
        RECT  0.830 2.180 1.050 2.820 ;
        RECT  1.050 2.220 1.660 2.820 ;
        RECT  1.660 2.030 1.880 2.820 ;
        RECT  1.880 2.220 2.490 2.820 ;
        RECT  2.490 2.030 2.710 2.820 ;
        RECT  2.710 2.220 4.220 2.820 ;
        RECT  4.220 2.030 4.440 2.820 ;
        RECT  4.440 2.220 5.020 2.820 ;
        RECT  5.020 2.180 5.240 2.820 ;
        RECT  5.240 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.900 0.660 4.020 1.560 ;
        RECT  4.020 1.420 4.150 1.560 ;
        RECT  1.320 0.450 1.420 0.870 ;
        RECT  1.420 0.450 1.540 1.640 ;
        RECT  1.540 1.080 2.410 1.240 ;
        RECT  1.540 0.470 3.420 0.590 ;
        RECT  3.420 0.470 3.540 1.380 ;
        RECT  3.540 1.260 3.600 1.380 ;
        RECT  3.540 0.630 3.710 0.790 ;
        RECT  3.600 1.260 3.760 1.570 ;
        RECT  2.020 0.720 2.710 0.880 ;
        RECT  2.710 0.720 2.870 1.560 ;
        RECT  2.870 1.400 2.990 1.560 ;
        RECT  3.850 0.660 3.900 1.140 ;
        RECT  4.840 1.760 5.510 1.920 ;
        RECT  4.740 0.710 5.500 0.870 ;
        RECT  4.740 1.500 4.840 1.920 ;
        RECT  6.120 0.680 6.270 0.840 ;
        RECT  6.120 1.390 6.220 1.810 ;
        RECT  6.060 0.470 6.120 1.810 ;
        RECT  6.000 0.470 6.060 1.510 ;
        RECT  4.390 0.470 6.000 0.590 ;
        RECT  4.270 0.470 4.390 1.810 ;
        RECT  3.400 1.690 4.270 1.810 ;
        RECT  3.300 1.640 3.400 1.810 ;
        RECT  3.180 0.710 3.300 1.810 ;
        RECT  6.400 0.630 6.560 1.720 ;
        RECT  6.930 1.050 7.010 1.270 ;
        RECT  6.790 1.050 6.930 2.050 ;
        RECT  5.840 1.930 6.790 2.050 ;
        RECT  5.760 0.710 5.870 0.870 ;
        RECT  5.760 1.610 5.840 2.050 ;
        RECT  5.680 0.710 5.760 2.050 ;
        RECT  6.240 1.090 6.400 1.250 ;
        RECT  3.060 0.710 3.180 0.870 ;
        RECT  4.620 0.710 4.740 1.920 ;
        RECT  3.680 0.980 3.850 1.140 ;
        RECT  5.640 0.710 5.680 1.730 ;
        RECT  1.250 1.490 1.420 1.640 ;
        RECT  2.030 1.400 2.710 1.560 ;
    END
END HCOSCOND1

MACRO HCOSCOND2
    CLASS CORE ;
    FOREIGN HCOSCOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.620 1.940 7.650 2.100 ;
        RECT  7.650 1.390 7.770 2.100 ;
        RECT  7.650 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.810 2.100 ;
        RECT  7.810 1.940 7.840 2.100 ;
        RECT  7.810 0.780 7.910 1.520 ;
        END
    END S
    PIN CS
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.670 1.515 ;
        RECT  5.670 1.145 5.960 1.305 ;
        END
    END CS
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.430 1.530 ;
        RECT  0.430 0.725 0.550 1.810 ;
        RECT  0.550 1.410 0.650 1.810 ;
        RECT  0.550 0.725 0.680 0.870 ;
        RECT  0.680 0.450 0.900 0.870 ;
        RECT  0.650 1.410 1.120 1.530 ;
        RECT  1.120 1.410 1.340 1.810 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 2.050 ;
        RECT  0.250 1.930 1.460 2.050 ;
        RECT  1.390 1.050 1.460 1.270 ;
        RECT  1.460 1.050 1.580 2.050 ;
        RECT  1.580 1.930 1.890 2.050 ;
        RECT  1.890 1.760 2.010 2.050 ;
        RECT  2.010 1.760 3.400 1.880 ;
        RECT  3.400 1.760 3.520 2.050 ;
        RECT  3.520 1.930 4.410 2.050 ;
        RECT  4.410 1.930 4.630 2.070 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.050 1.240 ;
        RECT  1.050 0.755 1.190 1.240 ;
        RECT  1.190 0.755 1.780 0.875 ;
        RECT  1.780 0.755 1.940 1.290 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.770 0.300 ;
        RECT  4.770 -0.300 4.990 0.340 ;
        RECT  4.990 -0.300 5.560 0.300 ;
        RECT  5.560 -0.300 5.780 0.340 ;
        RECT  5.780 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.200 2.820 ;
        RECT  2.200 2.030 2.420 2.820 ;
        RECT  2.420 2.220 3.030 2.820 ;
        RECT  3.030 2.030 3.250 2.820 ;
        RECT  3.250 2.220 4.760 2.820 ;
        RECT  4.760 2.030 4.980 2.820 ;
        RECT  4.980 2.220 5.560 2.820 ;
        RECT  5.560 2.180 5.780 2.820 ;
        RECT  5.780 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.660 1.390 6.760 1.810 ;
        RECT  6.660 0.675 6.810 0.835 ;
        RECT  5.280 1.500 5.380 1.920 ;
        RECT  5.280 0.710 6.040 0.870 ;
        RECT  5.380 1.760 6.050 1.920 ;
        RECT  4.390 0.660 4.440 1.140 ;
        RECT  4.440 0.660 4.560 1.560 ;
        RECT  4.560 1.420 4.690 1.560 ;
        RECT  1.840 0.470 2.170 0.630 ;
        RECT  2.170 0.470 2.290 1.640 ;
        RECT  2.290 1.080 2.950 1.240 ;
        RECT  2.290 0.470 3.960 0.590 ;
        RECT  3.960 0.470 4.080 1.380 ;
        RECT  4.080 1.260 4.140 1.380 ;
        RECT  4.080 0.630 4.250 0.790 ;
        RECT  4.140 1.260 4.300 1.570 ;
        RECT  2.560 0.720 3.250 0.880 ;
        RECT  3.250 0.720 3.410 1.560 ;
        RECT  3.410 1.400 3.530 1.560 ;
        RECT  6.600 0.470 6.660 1.810 ;
        RECT  6.540 0.470 6.600 1.510 ;
        RECT  4.930 0.470 6.540 0.590 ;
        RECT  4.810 0.470 4.930 1.810 ;
        RECT  3.970 1.690 4.810 1.810 ;
        RECT  3.840 1.640 3.970 1.810 ;
        RECT  3.720 0.710 3.840 1.810 ;
        RECT  6.940 0.625 7.100 1.720 ;
        RECT  7.470 1.050 7.550 1.270 ;
        RECT  7.330 1.050 7.470 2.050 ;
        RECT  6.380 1.930 7.330 2.050 ;
        RECT  6.300 0.710 6.410 0.870 ;
        RECT  6.300 1.610 6.380 2.050 ;
        RECT  6.220 0.710 6.300 2.050 ;
        RECT  6.180 0.710 6.220 1.730 ;
        RECT  6.780 1.090 6.940 1.250 ;
        RECT  3.600 0.710 3.720 0.870 ;
        RECT  5.160 0.710 5.280 1.920 ;
        RECT  4.220 0.980 4.390 1.140 ;
        RECT  1.790 1.480 2.170 1.640 ;
        RECT  2.570 1.400 3.250 1.560 ;
    END
END HCOSCOND2

MACRO HICIND1
    CLASS CORE ;
    FOREIGN HICIND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.895 1.940 4.925 2.100 ;
        RECT  4.925 1.390 5.085 2.100 ;
        RECT  4.925 0.420 5.085 0.920 ;
        RECT  5.085 1.940 5.115 2.100 ;
        RECT  5.085 1.390 5.210 1.515 ;
        RECT  5.085 0.800 5.210 0.920 ;
        RECT  5.210 0.800 5.350 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.060 1.940 0.090 2.100 ;
        RECT  0.060 0.420 0.090 1.510 ;
        RECT  0.090 0.420 0.180 2.100 ;
        RECT  0.180 1.390 0.250 2.100 ;
        RECT  0.180 0.420 0.250 0.640 ;
        RECT  0.250 1.940 0.285 2.100 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.130 1.515 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.235 2.820 ;
        RECT  1.235 2.180 1.455 2.820 ;
        RECT  1.455 2.220 2.810 2.820 ;
        RECT  2.810 2.180 3.030 2.820 ;
        RECT  3.030 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 0.710 3.270 0.870 ;
        RECT  2.750 1.650 3.280 1.810 ;
        RECT  0.835 1.460 0.975 1.700 ;
        RECT  0.975 1.460 1.075 1.580 ;
        RECT  0.440 0.760 1.075 0.880 ;
        RECT  1.075 0.440 1.195 1.580 ;
        RECT  1.195 0.440 1.295 0.880 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.390 0.710 2.630 0.870 ;
        RECT  3.620 1.930 3.860 2.090 ;
        RECT  0.715 1.930 3.620 2.050 ;
        RECT  0.715 1.065 0.845 1.225 ;
        RECT  3.930 0.470 4.010 0.690 ;
        RECT  3.930 1.350 4.000 1.570 ;
        RECT  3.810 0.470 3.930 1.570 ;
        RECT  1.935 0.470 3.810 0.590 ;
        RECT  1.935 1.080 2.445 1.240 ;
        RECT  1.815 0.470 1.935 1.810 ;
        RECT  1.715 0.470 1.815 0.910 ;
        RECT  4.250 0.470 4.420 0.630 ;
        RECT  4.250 1.410 4.410 1.570 ;
        RECT  4.130 0.470 4.250 1.570 ;
        RECT  4.675 1.080 4.890 1.240 ;
        RECT  4.555 1.080 4.675 1.810 ;
        RECT  3.660 1.690 4.555 1.810 ;
        RECT  3.540 0.720 3.690 0.880 ;
        RECT  3.540 1.650 3.660 1.810 ;
        RECT  4.070 1.015 4.130 1.235 ;
        RECT  1.615 1.650 1.815 1.810 ;
        RECT  0.595 1.065 0.715 2.050 ;
        RECT  2.390 1.650 2.630 1.810 ;
        RECT  0.300 0.760 0.440 1.275 ;
        RECT  3.400 0.720 3.540 1.810 ;
    END
END HICIND1

MACRO HICIND2
    CLASS CORE ;
    FOREIGN HICIND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.940 5.340 2.100 ;
        RECT  5.340 1.390 5.500 2.100 ;
        RECT  5.340 0.420 5.500 0.900 ;
        RECT  5.500 1.940 5.530 2.100 ;
        RECT  5.500 1.390 5.530 1.515 ;
        RECT  5.500 0.780 5.530 0.900 ;
        RECT  5.530 0.780 5.670 1.515 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.940 0.450 2.100 ;
        RECT  0.410 0.750 0.450 1.515 ;
        RECT  0.450 0.750 0.550 2.100 ;
        RECT  0.550 1.390 0.610 2.100 ;
        RECT  0.610 1.940 0.640 2.100 ;
        RECT  0.550 0.750 0.660 0.910 ;
        END
    END CO
    PIN CIN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        RECT  3.430 1.035 3.490 1.255 ;
        END
    END CIN
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.730 0.300 ;
        RECT  5.730 -0.300 5.950 0.340 ;
        RECT  5.950 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.545 2.820 ;
        RECT  1.545 2.180 1.765 2.820 ;
        RECT  1.765 2.220 3.170 2.820 ;
        RECT  3.170 2.180 3.390 2.820 ;
        RECT  3.390 2.220 4.920 2.820 ;
        RECT  4.920 2.180 5.140 2.820 ;
        RECT  5.140 2.220 5.730 2.820 ;
        RECT  5.730 2.180 5.950 2.820 ;
        RECT  5.950 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.555 0.440 1.655 0.880 ;
        RECT  1.435 0.440 1.555 1.580 ;
        RECT  0.290 0.470 1.435 0.590 ;
        RECT  1.335 1.460 1.435 1.580 ;
        RECT  1.175 1.460 1.335 1.700 ;
        RECT  3.110 1.650 3.660 1.810 ;
        RECT  3.110 0.710 3.650 0.870 ;
        RECT  2.990 0.710 3.110 1.810 ;
        RECT  2.750 0.710 2.990 0.870 ;
        RECT  3.980 1.930 4.220 2.090 ;
        RECT  1.055 1.930 3.980 2.050 ;
        RECT  1.055 1.065 1.205 1.225 ;
        RECT  4.340 0.470 4.390 0.690 ;
        RECT  4.340 1.350 4.380 1.570 ;
        RECT  4.220 0.470 4.340 1.570 ;
        RECT  2.295 0.470 4.220 0.590 ;
        RECT  2.295 1.080 2.855 1.240 ;
        RECT  2.175 0.440 2.295 1.810 ;
        RECT  2.075 0.440 2.175 0.880 ;
        RECT  4.650 0.470 4.780 0.630 ;
        RECT  4.650 1.410 4.770 1.570 ;
        RECT  4.530 0.470 4.650 1.570 ;
        RECT  5.035 1.080 5.400 1.240 ;
        RECT  4.915 1.080 5.035 1.810 ;
        RECT  4.020 1.690 4.915 1.810 ;
        RECT  3.940 0.720 4.050 0.880 ;
        RECT  3.940 1.650 4.020 1.810 ;
        RECT  4.480 1.015 4.530 1.235 ;
        RECT  1.975 1.650 2.175 1.810 ;
        RECT  0.935 1.065 1.055 2.050 ;
        RECT  2.750 1.650 2.990 1.810 ;
        RECT  0.140 0.470 0.290 1.275 ;
        RECT  3.800 0.720 3.940 1.810 ;
    END
END HICIND2

MACRO HICOND1
    CLASS CORE ;
    FOREIGN HICOND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.940 4.550 2.100 ;
        RECT  4.550 0.420 4.710 2.100 ;
        RECT  4.710 1.940 4.740 2.100 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.780 0.170 1.525 ;
        RECT  0.170 0.420 0.230 1.525 ;
        RECT  0.230 0.420 0.330 0.900 ;
        RECT  0.560 1.940 0.590 2.100 ;
        RECT  0.230 1.390 0.590 1.525 ;
        RECT  0.590 1.390 0.750 2.100 ;
        RECT  0.750 1.940 0.780 2.100 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.740 1.050 0.940 1.270 ;
        RECT  0.940 1.050 1.050 2.050 ;
        RECT  1.050 1.005 1.060 2.050 ;
        RECT  1.060 1.005 1.190 1.515 ;
        RECT  1.060 1.930 3.530 2.050 ;
        RECT  3.530 1.930 3.770 2.090 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.500 1.270 ;
        RECT  0.500 0.750 0.620 1.270 ;
        RECT  0.620 0.750 1.360 0.870 ;
        RECT  1.360 0.750 1.520 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.840 0.300 ;
        RECT  0.840 -0.300 1.060 0.340 ;
        RECT  1.060 -0.300 2.340 0.300 ;
        RECT  2.340 -0.300 2.560 0.340 ;
        RECT  2.560 -0.300 4.115 0.300 ;
        RECT  4.115 -0.300 4.335 0.340 ;
        RECT  4.335 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 4.115 2.820 ;
        RECT  4.115 2.180 4.335 2.820 ;
        RECT  4.335 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.065 1.050 4.185 1.810 ;
        RECT  4.185 1.050 4.430 1.270 ;
        RECT  3.710 0.490 3.830 1.570 ;
        RECT  3.830 1.410 3.930 1.570 ;
        RECT  3.830 0.490 3.930 0.910 ;
        RECT  1.230 1.650 1.685 1.810 ;
        RECT  1.470 0.470 1.685 0.590 ;
        RECT  1.685 0.470 1.805 1.810 ;
        RECT  1.805 1.080 2.290 1.240 ;
        RECT  1.805 0.470 3.350 0.590 ;
        RECT  3.350 0.470 3.470 1.570 ;
        RECT  3.470 1.410 3.580 1.570 ;
        RECT  3.470 0.660 3.590 0.820 ;
        RECT  1.940 0.720 2.610 0.880 ;
        RECT  2.610 0.720 2.770 1.790 ;
        RECT  3.190 1.690 4.065 1.810 ;
        RECT  3.090 0.720 3.210 0.860 ;
        RECT  3.090 1.650 3.190 1.810 ;
        RECT  2.970 0.720 3.090 1.810 ;
        RECT  3.600 1.090 3.710 1.250 ;
        RECT  1.230 0.440 1.470 0.590 ;
        RECT  1.940 1.630 2.610 1.790 ;
    END
END HICOND1

MACRO HICOND2
    CLASS CORE ;
    FOREIGN HICOND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.950 1.940 4.980 2.100 ;
        RECT  4.980 1.390 5.140 2.100 ;
        RECT  4.980 0.420 5.140 0.900 ;
        RECT  5.140 1.940 5.170 2.100 ;
        RECT  5.140 1.390 5.210 1.515 ;
        RECT  5.140 0.780 5.210 0.900 ;
        RECT  5.210 0.780 5.350 1.515 ;
        END
    END S
    PIN CON
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.770 0.550 1.765 ;
        RECT  0.550 0.770 0.805 0.900 ;
        RECT  0.805 0.420 0.965 0.900 ;
        RECT  0.550 1.595 1.350 1.765 ;
        END
    END CON
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.245 2.050 ;
        RECT  0.245 1.930 1.480 2.050 ;
        RECT  1.360 1.045 1.480 1.265 ;
        RECT  1.480 1.045 1.620 2.050 ;
        RECT  1.620 1.930 4.080 2.050 ;
        RECT  4.080 1.930 4.320 2.090 ;
        END
    END CI
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.825 1.075 1.120 1.235 ;
        RECT  1.120 0.750 1.240 1.235 ;
        RECT  1.240 0.750 1.980 0.870 ;
        RECT  1.980 0.750 2.150 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.340 ;
        RECT  3.110 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.160 0.720 3.320 1.790 ;
        RECT  2.680 0.720 3.160 0.840 ;
        RECT  2.680 1.670 3.160 1.790 ;
        RECT  2.520 0.720 2.680 0.940 ;
        RECT  4.020 0.660 4.140 0.820 ;
        RECT  4.020 1.410 4.130 1.570 ;
        RECT  3.900 0.470 4.020 1.570 ;
        RECT  2.395 0.470 3.900 0.590 ;
        RECT  2.395 1.075 2.775 1.235 ;
        RECT  2.275 0.470 2.395 1.810 ;
        RECT  2.020 0.470 2.275 0.600 ;
        RECT  1.780 1.650 2.275 1.810 ;
        RECT  4.380 0.470 4.480 0.910 ;
        RECT  4.380 1.410 4.480 1.570 ;
        RECT  4.260 0.470 4.380 1.570 ;
        RECT  4.735 1.080 5.040 1.240 ;
        RECT  4.615 1.080 4.735 1.810 ;
        RECT  3.740 1.690 4.615 1.810 ;
        RECT  3.640 0.720 3.760 0.860 ;
        RECT  3.640 1.650 3.740 1.810 ;
        RECT  3.520 0.720 3.640 1.810 ;
        RECT  4.150 1.090 4.260 1.250 ;
        RECT  1.780 0.440 2.020 0.600 ;
        RECT  2.520 1.550 2.680 1.790 ;
    END
END HICOND2

MACRO IAO21D0
    CLASS CORE ;
    FOREIGN IAO21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.820 1.690 1.980 ;
        RECT  1.250 0.470 1.690 0.630 ;
        RECT  1.690 0.470 1.830 1.980 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.535 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.535 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.295 0.410 1.515 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.820 2.820 ;
        RECT  0.820 2.180 1.040 2.820 ;
        RECT  1.040 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.130 0.965 1.150 1.130 ;
        RECT  0.990 0.520 1.130 2.050 ;
        RECT  0.460 0.520 0.990 0.680 ;
        RECT  0.130 1.890 0.990 2.050 ;
    END
END IAO21D0

MACRO IAO21D1
    CLASS CORE ;
    FOREIGN IAO21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.420 1.450 0.845 ;
        RECT  1.480 1.635 1.690 2.055 ;
        RECT  1.450 0.725 1.690 0.845 ;
        RECT  1.690 0.725 1.700 2.055 ;
        RECT  1.700 0.725 1.830 1.755 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.370 0.730 1.610 ;
        RECT  0.730 1.005 0.870 1.610 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.295 0.410 1.515 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.820 2.820 ;
        RECT  0.820 2.180 1.040 2.820 ;
        RECT  1.040 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.110 1.050 1.150 2.015 ;
        RECT  0.990 0.470 1.110 2.015 ;
        RECT  0.460 0.470 0.990 0.630 ;
        RECT  0.130 1.855 0.990 2.015 ;
    END
END IAO21D1

MACRO IAO21D2
    CLASS CORE ;
    FOREIGN IAO21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 0.420 1.450 0.845 ;
        RECT  1.485 1.650 1.690 1.810 ;
        RECT  1.450 0.725 1.690 0.845 ;
        RECT  1.690 0.725 1.830 1.810 ;
        RECT  1.830 0.725 1.920 0.845 ;
        RECT  1.920 0.420 2.150 0.845 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.370 0.730 1.610 ;
        RECT  0.730 1.005 0.870 1.610 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.295 0.410 1.515 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.820 2.820 ;
        RECT  0.820 2.180 1.040 2.820 ;
        RECT  1.040 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.040 1.030 2.200 2.050 ;
        RECT  1.150 1.930 2.040 2.050 ;
        RECT  1.110 1.050 1.150 2.050 ;
        RECT  0.990 0.470 1.110 2.050 ;
        RECT  0.460 0.470 0.990 0.630 ;
        RECT  0.130 1.855 0.990 2.015 ;
    END
END IAO21D2

MACRO IAO21D4
    CLASS CORE ;
    FOREIGN IAO21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.900 0.710 2.190 0.870 ;
        RECT  2.190 0.710 2.270 1.770 ;
        RECT  2.270 0.710 2.330 2.070 ;
        RECT  2.330 1.650 2.490 2.070 ;
        RECT  2.330 0.710 2.840 0.870 ;
        RECT  2.490 1.650 3.600 1.770 ;
        RECT  3.600 1.650 3.820 2.070 ;
        RECT  3.820 1.650 4.110 1.935 ;
        RECT  3.270 0.710 4.110 0.870 ;
        RECT  4.110 0.710 4.270 1.935 ;
        RECT  4.270 1.425 4.530 1.935 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.460 1.050 2.650 1.270 ;
        RECT  2.650 1.005 2.790 1.515 ;
        RECT  2.790 1.395 3.480 1.515 ;
        RECT  3.480 1.030 3.640 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 0.840 0.410 1.000 ;
        RECT  0.410 0.840 0.550 1.515 ;
        RECT  0.550 0.840 1.520 1.000 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.285 0.920 1.515 ;
        RECT  0.920 1.240 1.080 1.515 ;
        RECT  1.080 1.285 1.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.125 0.300 ;
        RECT  0.125 -0.300 0.345 0.340 ;
        RECT  0.345 -0.300 4.430 0.300 ;
        RECT  4.430 -0.300 4.650 0.340 ;
        RECT  4.650 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.290 2.820 ;
        RECT  0.290 2.180 0.510 2.820 ;
        RECT  0.510 2.220 1.610 2.820 ;
        RECT  1.610 2.180 1.830 2.820 ;
        RECT  1.830 2.220 2.940 2.820 ;
        RECT  2.940 2.180 3.160 2.820 ;
        RECT  3.160 2.220 4.260 2.820 ;
        RECT  4.260 2.180 4.480 2.820 ;
        RECT  4.480 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.390 0.470 4.550 1.230 ;
        RECT  3.130 0.470 4.390 0.590 ;
        RECT  2.970 0.470 3.130 1.270 ;
        RECT  1.770 0.470 2.970 0.590 ;
        RECT  1.770 1.080 2.000 1.240 ;
        RECT  1.650 0.470 1.770 1.755 ;
        RECT  0.500 0.510 1.650 0.670 ;
        RECT  1.160 1.635 1.650 1.755 ;
        RECT  0.940 1.635 1.160 2.055 ;
        LAYER M1 ;
        RECT  4.110 0.710 4.270 1.255 ;
        RECT  3.820 1.650 3.895 1.935 ;
        RECT  3.600 1.650 3.820 2.070 ;
        RECT  2.490 1.650 3.600 1.770 ;
        RECT  2.330 0.710 2.840 0.870 ;
        RECT  2.330 1.650 2.490 2.070 ;
        RECT  2.270 0.710 2.330 2.070 ;
        RECT  2.190 0.710 2.270 1.770 ;
        RECT  1.900 0.710 2.190 0.870 ;
        RECT  3.270 0.710 4.110 0.870 ;
    END
END IAO21D4

MACRO IAO22D0
    CLASS CORE ;
    FOREIGN IAO22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.950 1.600 1.370 1.760 ;
        RECT  1.250 0.420 1.370 0.580 ;
        RECT  1.370 0.420 1.510 1.760 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.985 2.150 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.950 1.690 1.170 ;
        RECT  1.690 0.725 1.830 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.985 0.570 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.535 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.720 2.820 ;
        RECT  0.720 2.180 0.940 2.820 ;
        RECT  0.940 2.220 1.660 2.820 ;
        RECT  1.660 1.600 1.880 2.820 ;
        RECT  1.880 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.810 1.080 1.250 1.240 ;
        RECT  0.690 0.450 0.810 2.050 ;
        RECT  0.480 0.450 0.690 0.610 ;
        RECT  0.070 1.890 0.690 2.050 ;
    END
END IAO22D0

MACRO IAO22D1
    CLASS CORE ;
    FOREIGN IAO22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.960 1.090 2.100 ;
        RECT  1.090 1.390 1.250 2.100 ;
        RECT  1.250 1.960 1.280 2.100 ;
        RECT  1.250 1.390 1.370 1.515 ;
        RECT  1.370 0.750 1.470 1.515 ;
        RECT  1.470 0.450 1.510 1.515 ;
        RECT  1.510 0.450 1.700 0.870 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        RECT  0.960 -0.300 1.180 0.340 ;
        RECT  1.180 -0.300 2.140 0.300 ;
        RECT  2.140 -0.300 2.360 0.340 ;
        RECT  2.360 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.700 2.820 ;
        RECT  0.700 2.180 0.920 2.820 ;
        RECT  0.920 2.220 1.850 2.820 ;
        RECT  1.850 2.180 2.070 2.820 ;
        RECT  2.070 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.060 0.495 1.220 1.270 ;
        RECT  0.560 0.495 1.060 0.655 ;
        RECT  0.440 0.495 0.560 1.640 ;
        RECT  0.280 1.520 0.440 1.640 ;
        RECT  2.460 1.960 2.490 2.100 ;
        RECT  2.300 1.370 2.460 2.100 ;
        RECT  1.660 1.635 2.300 1.755 ;
        RECT  2.270 1.960 2.300 2.100 ;
        RECT  0.060 1.520 0.280 1.940 ;
        RECT  1.440 1.635 1.660 2.055 ;
    END
END IAO22D1

MACRO IAO22D2
    CLASS CORE ;
    FOREIGN IAO22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.960 2.590 2.100 ;
        RECT  2.590 1.390 2.650 2.100 ;
        RECT  2.610 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.750 2.100 ;
        RECT  2.750 1.960 2.780 2.100 ;
        RECT  2.750 0.780 2.790 1.515 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.005 2.140 1.515 ;
        RECT  2.140 1.050 2.190 1.270 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.340 ;
        RECT  2.390 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.370 2.820 ;
        RECT  1.370 2.180 1.590 2.820 ;
        RECT  1.590 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.820 0.470 0.980 0.690 ;
        RECT  0.260 0.470 0.820 0.590 ;
        RECT  1.490 1.640 2.020 1.800 ;
        RECT  1.490 0.710 1.770 0.870 ;
        RECT  1.370 0.710 1.490 1.800 ;
        RECT  2.490 1.080 2.510 1.240 ;
        RECT  2.350 0.470 2.490 1.290 ;
        RECT  1.390 0.470 2.350 0.590 ;
        RECT  1.220 0.430 1.390 0.590 ;
        RECT  1.150 0.430 1.220 0.930 ;
        RECT  1.150 1.960 1.180 2.100 ;
        RECT  1.100 0.430 1.150 2.100 ;
        RECT  0.990 0.810 1.100 2.100 ;
        RECT  0.960 1.960 0.990 2.100 ;
        RECT  1.270 1.080 1.370 1.240 ;
        RECT  0.100 0.470 0.260 0.950 ;
    END
END IAO22D2

MACRO IAO22D4
    CLASS CORE ;
    FOREIGN IAO22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 1.640 4.110 2.020 ;
        RECT  3.625 0.500 4.110 0.880 ;
        RECT  4.110 0.500 4.530 2.020 ;
        RECT  4.530 1.640 4.590 2.020 ;
        RECT  4.530 0.500 4.600 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.005 2.800 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.110 1.515 ;
        RECT  3.110 1.050 3.245 1.270 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        RECT  0.240 1.395 1.265 1.515 ;
        RECT  1.265 1.030 1.425 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.225 0.300 ;
        RECT  3.225 -0.300 3.445 0.340 ;
        RECT  3.445 -0.300 4.770 0.300 ;
        RECT  4.770 -0.300 4.990 0.340 ;
        RECT  4.990 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.225 2.820 ;
        RECT  3.225 2.180 3.445 2.820 ;
        RECT  3.445 2.220 4.770 2.820 ;
        RECT  4.770 2.180 4.990 2.820 ;
        RECT  4.990 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 0.470 2.455 0.590 ;
        RECT  0.765 0.470 0.985 0.850 ;
        RECT  0.290 0.470 0.765 0.590 ;
        RECT  2.325 1.640 3.110 1.800 ;
        RECT  2.325 0.710 2.815 0.870 ;
        RECT  2.205 0.710 2.325 1.800 ;
        RECT  3.505 1.080 3.715 1.240 ;
        RECT  3.385 1.080 3.505 2.040 ;
        RECT  1.740 1.920 3.385 2.040 ;
        RECT  1.710 0.710 2.075 0.870 ;
        RECT  1.710 1.920 1.740 2.100 ;
        RECT  1.550 0.710 1.710 2.100 ;
        RECT  1.520 1.930 1.550 2.100 ;
        RECT  0.290 1.930 1.520 2.050 ;
        RECT  1.880 1.080 2.205 1.240 ;
        RECT  0.070 0.470 0.290 0.850 ;
        RECT  0.430 1.650 1.380 1.810 ;
        RECT  0.070 1.650 0.290 2.050 ;
        LAYER M1 ;
        RECT  3.625 0.500 3.895 0.880 ;
        RECT  3.625 1.640 3.885 2.020 ;
    END
END IAO22D4

MACRO IIND4D0
    CLASS CORE ;
    FOREIGN IIND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.470 0.870 2.050 ;
        RECT  0.870 0.470 1.000 0.630 ;
        RECT  0.870 1.890 1.810 2.050 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.000 1.200 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.535 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.540 ;
        RECT  1.510 1.370 1.610 1.540 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.610 0.610 2.050 ;
        RECT  2.140 0.470 2.490 0.630 ;
        RECT  2.140 1.890 2.490 2.050 ;
        RECT  2.020 0.470 2.140 2.050 ;
        RECT  0.070 1.890 0.450 2.050 ;
        RECT  1.720 1.080 2.020 1.240 ;
    END
END IIND4D0

MACRO IIND4D1
    CLASS CORE ;
    FOREIGN IIND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.420 0.730 0.870 ;
        RECT  0.730 0.420 0.870 1.770 ;
        RECT  0.870 0.420 0.930 0.870 ;
        RECT  0.870 1.640 1.090 2.080 ;
        RECT  1.090 1.640 1.580 1.760 ;
        RECT  1.580 1.640 1.800 2.080 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.990 0.250 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.210 1.650 1.380 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.860 0.300 ;
        RECT  1.860 -0.300 2.080 0.340 ;
        RECT  2.080 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.550 1.200 0.610 1.420 ;
        RECT  0.430 0.660 0.550 2.050 ;
        RECT  0.390 0.660 0.430 0.900 ;
        RECT  2.140 0.470 2.490 0.630 ;
        RECT  2.140 1.890 2.490 2.050 ;
        RECT  2.020 0.470 2.140 2.050 ;
        RECT  1.770 1.095 2.020 1.255 ;
        RECT  0.070 1.890 0.430 2.050 ;
    END
END IIND4D1

MACRO IIND4D2
    CLASS CORE ;
    FOREIGN IIND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.045 1.650 1.050 2.070 ;
        RECT  1.040 0.750 1.050 0.970 ;
        RECT  1.050 0.750 1.190 2.070 ;
        RECT  1.190 0.750 1.200 0.970 ;
        RECT  1.190 1.650 1.265 2.070 ;
        RECT  1.265 1.650 1.875 1.770 ;
        RECT  1.875 1.650 2.095 2.070 ;
        RECT  2.095 1.650 2.705 1.770 ;
        RECT  2.705 1.650 2.925 2.070 ;
        RECT  2.925 1.650 3.535 1.770 ;
        RECT  3.535 1.650 3.755 2.070 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.110 2.810 1.515 ;
        RECT  2.810 1.285 3.110 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.285 1.990 1.515 ;
        RECT  1.990 1.120 2.150 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.725 4.710 1.250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        RECT  0.640 2.180 0.860 2.820 ;
        RECT  0.860 2.220 1.460 2.820 ;
        RECT  1.460 2.180 1.680 2.820 ;
        RECT  1.680 2.220 2.290 2.820 ;
        RECT  2.290 2.180 2.510 2.820 ;
        RECT  2.510 2.220 3.120 2.820 ;
        RECT  3.120 2.180 3.340 2.820 ;
        RECT  3.340 2.220 3.950 2.820 ;
        RECT  3.950 2.180 4.170 2.820 ;
        RECT  4.170 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.160 0.925 1.320 ;
        RECT  0.420 0.420 0.540 1.750 ;
        RECT  0.070 0.420 0.420 0.580 ;
        RECT  1.610 0.500 2.370 0.660 ;
        RECT  1.390 0.500 1.610 0.930 ;
        RECT  0.820 0.500 1.390 0.620 ;
        RECT  3.990 0.500 4.150 1.020 ;
        RECT  3.490 0.500 3.990 0.620 ;
        RECT  3.270 0.500 3.490 0.920 ;
        RECT  4.390 0.420 4.740 0.580 ;
        RECT  4.390 1.590 4.605 1.750 ;
        RECT  4.270 0.420 4.390 1.750 ;
        RECT  3.710 1.160 4.270 1.320 ;
        RECT  2.510 0.500 3.270 0.660 ;
        RECT  1.750 0.780 3.130 0.940 ;
        RECT  0.660 0.500 0.820 1.020 ;
        RECT  0.195 1.590 0.420 1.750 ;
    END
END IIND4D2

MACRO IIND4D4
    CLASS CORE ;
    FOREIGN IIND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.620 1.870 2.000 ;
        RECT  1.430 0.760 1.870 0.920 ;
        RECT  1.870 0.760 2.290 2.000 ;
        RECT  2.290 0.760 2.450 0.920 ;
        RECT  2.290 1.620 7.330 2.000 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.410 1.005 8.570 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.920 2.820 ;
        RECT  0.920 2.180 1.140 2.820 ;
        RECT  1.140 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.570 2.820 ;
        RECT  2.570 2.180 2.790 2.820 ;
        RECT  2.790 2.220 3.400 2.820 ;
        RECT  3.400 2.180 3.620 2.820 ;
        RECT  3.620 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.060 2.820 ;
        RECT  5.060 2.180 5.280 2.820 ;
        RECT  5.280 2.220 5.880 2.820 ;
        RECT  5.880 2.180 6.100 2.820 ;
        RECT  6.100 2.220 6.700 2.820 ;
        RECT  6.700 2.180 6.920 2.820 ;
        RECT  6.920 2.220 7.520 2.820 ;
        RECT  7.520 2.180 7.740 2.820 ;
        RECT  7.740 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.690 1.080 1.580 1.240 ;
        RECT  0.690 1.960 0.720 2.100 ;
        RECT  0.610 1.080 0.690 2.100 ;
        RECT  0.530 0.420 0.610 2.100 ;
        RECT  0.450 0.420 0.530 1.240 ;
        RECT  2.810 0.470 4.330 0.630 ;
        RECT  2.590 0.470 2.810 0.910 ;
        RECT  1.290 0.470 2.590 0.630 ;
        RECT  7.350 0.470 7.570 0.890 ;
        RECT  6.880 0.470 7.350 0.590 ;
        RECT  6.660 0.470 6.880 0.890 ;
        RECT  6.190 0.470 6.660 0.590 ;
        RECT  5.970 0.470 6.190 0.890 ;
        RECT  8.120 0.420 8.190 1.240 ;
        RECT  8.120 1.960 8.150 2.100 ;
        RECT  8.030 0.420 8.120 2.100 ;
        RECT  7.960 1.080 8.030 2.100 ;
        RECT  6.540 1.080 7.960 1.240 ;
        RECT  7.930 1.960 7.960 2.100 ;
        RECT  4.450 0.470 5.970 0.630 ;
        RECT  2.950 0.750 5.830 0.885 ;
        RECT  1.070 0.470 1.290 0.910 ;
        RECT  0.500 1.960 0.530 2.100 ;
        LAYER M1 ;
        RECT  1.330 1.620 1.655 2.000 ;
        RECT  1.430 0.760 1.655 0.920 ;
        RECT  2.505 1.620 7.330 2.000 ;
    END
END IIND4D4

MACRO IINR4D0
    CLASS CORE ;
    FOREIGN IINR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.460 0.830 1.535 ;
        RECT  0.830 0.440 0.870 1.535 ;
        RECT  0.870 0.440 1.050 0.600 ;
        RECT  1.050 0.470 1.590 0.600 ;
        RECT  1.590 0.440 1.830 0.600 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.720 1.510 1.235 ;
        RECT  1.510 0.720 1.630 0.940 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.725 2.470 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.095 1.810 1.795 ;
        RECT  1.810 0.930 1.830 1.795 ;
        RECT  1.830 0.930 1.950 1.215 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.840 2.820 ;
        RECT  1.840 2.180 2.060 2.820 ;
        RECT  2.060 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.190 1.500 2.500 1.660 ;
        RECT  2.280 0.430 2.500 0.590 ;
        RECT  0.450 0.470 0.610 2.100 ;
        RECT  2.190 0.470 2.280 0.590 ;
        RECT  2.070 0.470 2.190 2.050 ;
        RECT  1.200 1.930 2.070 2.050 ;
        RECT  0.070 0.470 0.450 0.630 ;
        RECT  1.040 0.720 1.200 2.050 ;
    END
END IINR4D0

MACRO IINR4D1
    CLASS CORE ;
    FOREIGN IINR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.655 1.370 0.815 ;
        RECT  1.370 0.655 1.510 1.570 ;
        RECT  1.510 0.655 1.840 0.815 ;
        RECT  1.510 1.410 2.070 1.570 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.960 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.725 3.130 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.725 3.430 1.270 ;
        RECT  3.430 1.050 3.520 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.440 0.300 ;
        RECT  0.440 -0.300 0.660 0.690 ;
        RECT  0.660 -0.300 2.000 0.300 ;
        RECT  2.000 -0.300 2.220 0.815 ;
        RECT  2.220 -0.300 3.100 0.300 ;
        RECT  3.100 -0.300 3.320 0.340 ;
        RECT  3.320 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.230 2.820 ;
        RECT  3.230 2.180 3.450 2.820 ;
        RECT  3.450 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.480 1.930 2.720 2.100 ;
        RECT  0.290 1.930 2.480 2.050 ;
        RECT  2.800 1.410 3.070 1.570 ;
        RECT  2.800 0.420 2.920 0.580 ;
        RECT  2.680 0.420 2.800 1.570 ;
        RECT  3.640 0.660 3.760 1.810 ;
        RECT  3.590 0.660 3.640 0.900 ;
        RECT  3.590 1.470 3.640 1.810 ;
        RECT  2.315 1.690 3.590 1.810 ;
        RECT  2.195 1.080 2.315 1.810 ;
        RECT  2.470 1.045 2.680 1.205 ;
        RECT  0.070 1.930 0.290 2.090 ;
        RECT  1.800 1.080 2.195 1.240 ;
    END
END IINR4D1

MACRO IINR4D2
    CLASS CORE ;
    FOREIGN IINR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.380 1.230 1.810 ;
        RECT  1.230 1.380 1.690 1.500 ;
        RECT  1.690 0.485 1.770 1.500 ;
        RECT  1.770 0.485 1.830 1.810 ;
        RECT  1.830 1.350 1.990 1.810 ;
        RECT  1.830 0.485 6.080 0.645 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 0.725 7.590 1.250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.280 0.300 ;
        RECT  1.280 -0.300 1.500 0.340 ;
        RECT  1.500 -0.300 2.100 0.300 ;
        RECT  2.100 -0.300 2.320 0.340 ;
        RECT  2.320 -0.300 2.610 0.300 ;
        RECT  2.610 -0.300 2.830 0.340 ;
        RECT  2.830 -0.300 3.430 0.300 ;
        RECT  3.430 -0.300 3.650 0.340 ;
        RECT  3.650 -0.300 3.910 0.300 ;
        RECT  3.910 -0.300 4.130 0.340 ;
        RECT  4.130 -0.300 4.730 0.300 ;
        RECT  4.730 -0.300 4.950 0.340 ;
        RECT  4.950 -0.300 5.430 0.300 ;
        RECT  5.430 -0.300 5.650 0.340 ;
        RECT  5.650 -0.300 6.250 0.300 ;
        RECT  6.250 -0.300 6.470 0.340 ;
        RECT  6.470 -0.300 7.310 0.300 ;
        RECT  7.310 -0.300 7.530 0.340 ;
        RECT  7.530 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.590 0.420 0.750 1.200 ;
        RECT  0.750 1.040 1.540 1.200 ;
        RECT  0.540 1.040 0.590 1.200 ;
        RECT  0.400 1.040 0.540 1.645 ;
        RECT  0.250 1.505 0.400 1.645 ;
        RECT  3.670 1.890 3.890 2.050 ;
        RECT  3.130 1.930 3.670 2.050 ;
        RECT  2.910 1.630 3.130 2.050 ;
        RECT  2.370 1.930 2.910 2.050 ;
        RECT  2.340 1.930 2.370 2.100 ;
        RECT  2.180 1.370 2.340 2.100 ;
        RECT  2.150 1.930 2.180 2.100 ;
        RECT  1.610 1.930 2.150 2.050 ;
        RECT  1.390 1.630 1.610 2.050 ;
        RECT  0.820 1.930 1.390 2.050 ;
        RECT  5.080 1.380 5.300 1.810 ;
        RECT  4.540 1.380 5.080 1.500 ;
        RECT  4.440 1.380 4.540 1.810 ;
        RECT  4.320 1.220 4.440 1.810 ;
        RECT  3.510 1.220 4.320 1.340 ;
        RECT  3.390 1.220 3.510 1.810 ;
        RECT  3.290 1.380 3.390 1.810 ;
        RECT  2.750 1.380 3.290 1.500 ;
        RECT  6.870 1.380 7.030 2.050 ;
        RECT  6.370 1.890 6.870 2.050 ;
        RECT  6.340 1.890 6.370 2.100 ;
        RECT  6.180 1.370 6.340 2.100 ;
        RECT  6.150 1.930 6.180 2.100 ;
        RECT  5.680 1.930 6.150 2.050 ;
        RECT  5.650 1.930 5.680 2.100 ;
        RECT  5.490 1.370 5.650 2.100 ;
        RECT  5.460 1.930 5.490 2.100 ;
        RECT  4.920 1.930 5.460 2.050 ;
        RECT  4.700 1.630 4.920 2.050 ;
        RECT  4.130 1.930 4.700 2.050 ;
        RECT  4.010 1.460 4.130 2.050 ;
        RECT  7.430 1.525 7.590 2.070 ;
        RECT  7.290 1.525 7.430 1.665 ;
        RECT  7.150 1.070 7.290 1.665 ;
        RECT  7.090 1.070 7.150 1.200 ;
        RECT  6.930 0.420 7.090 1.200 ;
        RECT  3.270 0.765 6.930 0.885 ;
        RECT  3.150 0.765 3.270 1.200 ;
        RECT  3.970 1.460 4.010 1.680 ;
        RECT  2.530 1.380 2.750 1.810 ;
        RECT  2.470 1.040 3.150 1.200 ;
        RECT  0.660 1.380 0.820 2.050 ;
        RECT  0.090 1.505 0.250 2.070 ;
    END
END IINR4D2

MACRO IINR4D4
    CLASS CORE ;
    FOREIGN IINR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.780 1.360 8.910 1.780 ;
        RECT  2.190 0.470 8.910 0.590 ;
        RECT  8.910 0.470 9.000 1.780 ;
        RECT  9.000 0.470 9.330 1.480 ;
        RECT  9.330 1.360 9.540 1.480 ;
        RECT  9.540 1.360 9.760 1.780 ;
        RECT  9.330 0.470 9.920 0.610 ;
        RECT  9.760 1.360 10.300 1.480 ;
        RECT  10.300 1.360 10.520 1.780 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.725 2.790 0.955 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 0.725 5.350 0.955 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  11.910 1.005 12.070 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.820 0.300 ;
        RECT  0.820 -0.300 1.040 0.340 ;
        RECT  1.040 -0.300 1.800 0.300 ;
        RECT  1.800 -0.300 2.020 0.340 ;
        RECT  2.020 -0.300 2.630 0.300 ;
        RECT  2.630 -0.300 2.850 0.340 ;
        RECT  2.850 -0.300 3.460 0.300 ;
        RECT  3.460 -0.300 3.680 0.340 ;
        RECT  3.680 -0.300 4.290 0.300 ;
        RECT  4.290 -0.300 4.510 0.340 ;
        RECT  4.510 -0.300 5.120 0.300 ;
        RECT  5.120 -0.300 5.340 0.340 ;
        RECT  5.340 -0.300 6.780 0.300 ;
        RECT  6.780 -0.300 7.000 0.340 ;
        RECT  7.000 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.830 0.340 ;
        RECT  7.830 -0.300 8.440 0.300 ;
        RECT  8.440 -0.300 8.660 0.340 ;
        RECT  8.660 -0.300 9.260 0.300 ;
        RECT  9.260 -0.300 9.480 0.340 ;
        RECT  9.480 -0.300 10.090 0.300 ;
        RECT  10.090 -0.300 10.310 0.340 ;
        RECT  10.310 -0.300 11.110 0.300 ;
        RECT  11.110 -0.300 11.330 0.340 ;
        RECT  11.330 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.820 2.820 ;
        RECT  0.820 2.180 1.040 2.820 ;
        RECT  1.040 2.220 11.110 2.820 ;
        RECT  11.110 2.180 11.330 2.820 ;
        RECT  11.330 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.760 1.620 5.980 2.040 ;
        RECT  5.220 1.920 5.760 2.040 ;
        RECT  5.000 1.620 5.220 2.040 ;
        RECT  4.460 1.920 5.000 2.040 ;
        RECT  4.240 1.620 4.460 2.040 ;
        RECT  3.700 1.920 4.240 2.040 ;
        RECT  3.480 1.360 3.700 2.040 ;
        RECT  2.960 1.920 3.480 2.040 ;
        RECT  2.740 1.360 2.960 2.040 ;
        RECT  2.220 1.920 2.740 2.040 ;
        RECT  2.000 1.360 2.220 2.040 ;
        RECT  1.480 1.920 2.000 2.040 ;
        RECT  6.510 0.780 7.670 0.940 ;
        RECT  6.390 0.780 6.510 1.220 ;
        RECT  1.750 1.100 6.390 1.220 ;
        RECT  1.630 1.100 1.750 1.455 ;
        RECT  0.610 1.335 1.630 1.455 ;
        RECT  0.610 0.420 0.640 0.840 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 0.420 0.610 2.100 ;
        RECT  0.420 0.420 0.450 0.840 ;
        RECT  8.020 1.360 8.240 1.780 ;
        RECT  7.480 1.360 8.020 1.480 ;
        RECT  7.260 1.360 7.480 1.780 ;
        RECT  6.720 1.360 7.260 1.480 ;
        RECT  6.500 1.360 6.720 1.780 ;
        RECT  5.600 1.360 6.500 1.480 ;
        RECT  5.380 1.360 5.600 1.780 ;
        RECT  4.840 1.360 5.380 1.480 ;
        RECT  4.620 1.360 4.840 1.780 ;
        RECT  4.080 1.360 4.620 1.480 ;
        RECT  10.680 1.360 10.900 2.040 ;
        RECT  10.140 1.900 10.680 2.040 ;
        RECT  9.920 1.620 10.140 2.040 ;
        RECT  9.380 1.900 9.920 2.040 ;
        RECT  9.160 1.620 9.380 2.040 ;
        RECT  8.620 1.900 9.160 2.040 ;
        RECT  8.400 1.620 8.620 2.040 ;
        RECT  7.860 1.900 8.400 2.040 ;
        RECT  7.640 1.620 7.860 2.040 ;
        RECT  7.100 1.900 7.640 2.040 ;
        RECT  6.880 1.620 7.100 2.040 ;
        RECT  6.340 1.900 6.880 2.040 ;
        RECT  11.700 0.420 11.730 0.840 ;
        RECT  11.700 1.960 11.730 2.100 ;
        RECT  11.540 0.420 11.700 2.100 ;
        RECT  11.510 0.420 11.540 0.940 ;
        RECT  11.510 1.960 11.540 2.100 ;
        RECT  6.120 1.620 6.340 2.040 ;
        RECT  3.860 1.360 4.080 1.780 ;
        RECT  0.420 1.960 0.450 2.100 ;
        RECT  1.260 1.620 1.480 2.040 ;
        RECT  9.640 0.780 11.510 0.940 ;
        LAYER M1 ;
        RECT  10.300 1.360 10.520 1.780 ;
        RECT  9.760 1.360 10.300 1.480 ;
        RECT  2.190 0.470 8.695 0.590 ;
        RECT  9.545 0.470 9.920 0.610 ;
        RECT  9.545 1.360 9.760 1.780 ;
    END
END IINR4D4

MACRO IND2D0
    CLASS CORE ;
    FOREIGN IND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.840 1.890 1.370 2.050 ;
        RECT  1.130 0.470 1.370 0.630 ;
        RECT  1.370 0.470 1.510 2.050 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.910 1.240 ;
        RECT  0.420 0.470 0.540 2.050 ;
        RECT  0.070 0.470 0.420 0.630 ;
        RECT  0.070 1.890 0.420 2.050 ;
    END
END IND2D0

MACRO IND2D1
    CLASS CORE ;
    FOREIGN IND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.635 1.080 2.055 ;
        RECT  1.080 1.635 1.370 1.755 ;
        RECT  1.150 0.425 1.370 0.845 ;
        RECT  1.370 0.725 1.510 1.755 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.700 1.080 0.910 1.240 ;
        RECT  0.580 0.470 0.700 1.795 ;
        RECT  0.070 0.470 0.580 0.630 ;
        RECT  0.070 1.635 0.580 1.795 ;
    END
END IND2D1

MACRO IND2D2
    CLASS CORE ;
    FOREIGN IND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 1.630 0.990 2.050 ;
        RECT  1.130 0.440 1.370 0.600 ;
        RECT  0.990 1.630 1.530 1.750 ;
        RECT  1.530 1.630 1.750 2.050 ;
        RECT  1.750 1.630 2.010 1.750 ;
        RECT  1.370 0.480 2.010 0.600 ;
        RECT  2.010 0.480 2.150 1.750 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.270 ;
        RECT  0.870 0.725 1.690 0.845 ;
        RECT  1.690 0.725 1.850 1.290 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.370 2.820 ;
        RECT  0.370 2.180 0.590 2.820 ;
        RECT  0.590 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.370 0.480 0.490 1.670 ;
        RECT  0.490 1.390 1.190 1.510 ;
        RECT  1.190 1.030 1.350 1.510 ;
        RECT  0.290 0.480 0.370 0.600 ;
        RECT  0.070 1.510 0.370 1.670 ;
        RECT  0.070 0.440 0.290 0.600 ;
    END
END IND2D2

MACRO IND2D4
    CLASS CORE ;
    FOREIGN IND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  1.140 1.370 1.300 2.100 ;
        RECT  1.300 1.880 1.330 2.100 ;
        RECT  1.330 1.880 1.800 2.040 ;
        RECT  1.800 1.630 2.020 2.040 ;
        RECT  2.020 1.880 2.510 2.040 ;
        RECT  2.510 1.630 2.730 2.040 ;
        RECT  2.730 1.880 3.150 2.040 ;
        RECT  3.150 1.425 3.570 2.040 ;
        RECT  3.570 1.425 3.660 1.545 ;
        RECT  1.480 0.470 3.660 0.630 ;
        RECT  3.660 0.470 3.780 1.545 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.710 1.235 ;
        RECT  1.710 1.005 1.830 1.510 ;
        RECT  1.830 1.390 2.730 1.510 ;
        RECT  2.730 1.030 2.890 1.510 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.150 0.300 ;
        RECT  2.150 -0.300 2.370 0.340 ;
        RECT  2.370 -0.300 3.490 0.300 ;
        RECT  3.490 -0.300 3.710 0.340 ;
        RECT  3.710 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.370 0.765 3.530 1.255 ;
        RECT  2.340 0.765 3.370 0.885 ;
        RECT  2.180 0.765 2.340 1.270 ;
        RECT  1.200 0.765 2.180 0.885 ;
        RECT  1.080 0.765 1.200 1.240 ;
        RECT  0.835 1.080 1.080 1.240 ;
        RECT  0.715 0.765 0.835 1.755 ;
        RECT  0.710 0.765 0.715 0.885 ;
        RECT  0.640 1.635 0.715 1.755 ;
        RECT  0.490 0.465 0.710 0.885 ;
        RECT  0.420 1.635 0.640 2.055 ;
        LAYER M1 ;
        RECT  1.480 0.470 3.660 0.630 ;
        RECT  1.110 1.960 1.140 2.100 ;
        RECT  1.140 1.370 1.300 2.100 ;
        RECT  1.300 1.880 1.330 2.100 ;
        RECT  1.330 1.880 1.800 2.040 ;
        RECT  1.800 1.630 2.020 2.040 ;
        RECT  2.020 1.880 2.510 2.040 ;
        RECT  2.510 1.630 2.730 2.040 ;
        RECT  2.730 1.880 2.935 2.040 ;
        RECT  3.660 0.470 3.780 1.210 ;
    END
END IND2D4

MACRO IND3D0
    CLASS CORE ;
    FOREIGN IND3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.890 1.690 2.050 ;
        RECT  1.480 0.460 1.690 0.620 ;
        RECT  1.690 0.460 1.830 2.050 ;
        RECT  1.830 1.890 1.850 2.050 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.590 0.300 ;
        RECT  0.590 -0.300 0.810 0.340 ;
        RECT  0.810 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.240 2.820 ;
        RECT  1.240 2.180 1.460 2.820 ;
        RECT  1.460 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.880 1.240 ;
        RECT  0.420 0.460 0.540 2.050 ;
        RECT  0.150 0.460 0.420 0.620 ;
        RECT  0.070 1.890 0.420 2.050 ;
    END
END IND3D0

MACRO IND3D1
    CLASS CORE ;
    FOREIGN IND3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.850 1.960 0.880 2.100 ;
        RECT  0.880 1.390 1.040 2.100 ;
        RECT  1.040 1.960 1.070 2.100 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.040 1.390 1.670 1.510 ;
        RECT  1.670 1.390 1.690 2.100 ;
        RECT  1.660 0.420 1.690 0.900 ;
        RECT  1.690 0.420 1.830 2.100 ;
        RECT  1.830 1.960 1.860 2.100 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.725 1.530 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.725 1.210 1.270 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.240 2.820 ;
        RECT  1.240 2.180 1.460 2.820 ;
        RECT  1.460 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.730 1.080 0.880 1.240 ;
        RECT  0.610 0.470 0.730 1.660 ;
        RECT  0.290 0.470 0.610 0.605 ;
        RECT  0.070 1.500 0.610 1.660 ;
        RECT  0.070 0.445 0.290 0.605 ;
    END
END IND3D1

MACRO IND3D2
    CLASS CORE ;
    FOREIGN IND3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.670 1.020 2.090 ;
        RECT  1.020 1.670 1.530 1.790 ;
        RECT  1.530 1.670 1.750 2.090 ;
        RECT  1.510 0.430 1.750 0.590 ;
        RECT  1.750 1.670 2.230 1.790 ;
        RECT  2.230 1.670 2.450 2.090 ;
        RECT  2.450 1.670 2.650 1.790 ;
        RECT  1.750 0.470 2.650 0.590 ;
        RECT  2.650 0.470 2.790 1.790 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        RECT  1.200 1.395 2.030 1.515 ;
        RECT  2.030 1.030 2.190 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.255 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.730 0.340 ;
        RECT  0.730 -0.300 2.520 0.300 ;
        RECT  2.520 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.400 2.820 ;
        RECT  0.400 2.180 0.620 2.820 ;
        RECT  0.620 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.680 0.710 2.390 0.830 ;
        RECT  2.390 0.710 2.530 1.290 ;
        RECT  0.680 1.080 0.910 1.240 ;
        RECT  0.560 0.470 0.680 1.660 ;
        RECT  0.310 0.470 0.560 0.605 ;
        RECT  0.070 1.500 0.560 1.660 ;
        RECT  0.070 0.445 0.310 0.605 ;
    END
END IND3D2

MACRO IND3D4
    CLASS CORE ;
    FOREIGN IND3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.425 1.330 2.050 ;
        RECT  1.330 1.890 1.800 2.050 ;
        RECT  1.720 0.430 1.960 0.590 ;
        RECT  1.800 1.650 2.020 2.050 ;
        RECT  1.960 0.470 3.870 0.590 ;
        RECT  3.870 0.430 4.090 0.590 ;
        RECT  2.020 1.890 4.590 2.050 ;
        RECT  4.590 1.570 4.750 2.050 ;
        RECT  4.750 1.570 4.990 1.690 ;
        RECT  4.090 0.470 4.990 0.590 ;
        RECT  4.990 0.470 5.110 1.690 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.820 0.950 1.980 1.285 ;
        RECT  1.980 0.950 2.610 1.070 ;
        RECT  2.610 0.950 2.730 1.530 ;
        RECT  2.730 1.410 3.130 1.530 ;
        RECT  3.130 0.950 3.250 1.530 ;
        RECT  3.250 0.950 3.910 1.070 ;
        RECT  3.910 0.950 4.070 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.080 1.555 1.240 ;
        RECT  1.555 1.080 1.675 1.525 ;
        RECT  1.675 1.405 2.270 1.525 ;
        RECT  2.270 1.190 2.490 1.770 ;
        RECT  2.490 1.650 3.370 1.770 ;
        RECT  3.370 1.190 3.590 1.770 ;
        RECT  3.590 1.650 4.250 1.770 ;
        RECT  4.250 1.005 4.390 1.770 ;
        RECT  4.390 1.070 4.550 1.290 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.780 0.300 ;
        RECT  2.780 -0.300 3.000 0.340 ;
        RECT  3.000 -0.300 4.860 0.300 ;
        RECT  4.860 -0.300 5.080 0.340 ;
        RECT  5.080 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.965 2.820 ;
        RECT  4.965 2.180 5.200 2.820 ;
        RECT  5.200 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.850 0.710 3.010 1.285 ;
        RECT  3.010 0.710 4.710 0.830 ;
        RECT  4.710 0.710 4.870 1.305 ;
        RECT  1.120 0.710 2.850 0.830 ;
        RECT  1.000 0.710 1.120 1.240 ;
        RECT  0.620 1.080 1.000 1.240 ;
        RECT  0.610 0.420 0.620 1.240 ;
        RECT  0.460 0.420 0.610 2.055 ;
        RECT  0.450 1.080 0.460 2.055 ;
        LAYER M1 ;
        RECT  1.545 1.890 1.800 2.050 ;
        RECT  1.720 0.430 1.960 0.590 ;
        RECT  1.800 1.650 2.020 2.050 ;
        RECT  1.960 0.470 3.870 0.590 ;
        RECT  3.870 0.430 4.090 0.590 ;
        RECT  2.020 1.890 4.590 2.050 ;
        RECT  4.590 1.570 4.750 2.050 ;
        RECT  4.750 1.570 4.990 1.690 ;
        RECT  4.090 0.470 4.990 0.590 ;
        RECT  4.990 0.470 5.110 1.690 ;
    END
END IND3D4

MACRO IND4D0
    CLASS CORE ;
    FOREIGN IND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.890 2.010 2.050 ;
        RECT  1.810 0.470 2.010 0.630 ;
        RECT  2.010 0.470 2.150 2.050 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.550 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.600 0.300 ;
        RECT  0.600 -0.300 0.820 0.340 ;
        RECT  0.820 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.880 1.240 ;
        RECT  0.420 0.470 0.540 2.050 ;
        RECT  0.160 0.470 0.420 0.630 ;
        RECT  0.070 1.890 0.420 2.050 ;
    END
END IND4D0

MACRO IND4D1
    CLASS CORE ;
    FOREIGN IND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 1.635 1.030 2.050 ;
        RECT  1.030 1.635 1.550 1.755 ;
        RECT  1.550 1.635 1.770 2.050 ;
        RECT  1.770 1.635 2.010 1.755 ;
        RECT  1.850 0.420 2.010 0.840 ;
        RECT  2.010 0.420 2.070 1.755 ;
        RECT  2.070 0.720 2.150 1.755 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.890 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.550 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.900 1.240 ;
        RECT  0.420 0.710 0.540 1.800 ;
        RECT  0.070 0.710 0.420 0.870 ;
        RECT  0.070 1.640 0.420 1.800 ;
    END
END IND4D1

MACRO IND4D2
    CLASS CORE ;
    FOREIGN IND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.960 1.300 2.100 ;
        RECT  1.300 1.390 1.360 2.100 ;
        RECT  1.360 0.710 1.460 2.100 ;
        RECT  1.460 1.930 1.490 2.100 ;
        RECT  1.460 0.710 1.520 1.515 ;
        RECT  1.490 1.930 2.100 2.050 ;
        RECT  2.100 1.930 2.130 2.100 ;
        RECT  2.130 1.370 2.290 2.100 ;
        RECT  2.290 1.930 2.320 2.100 ;
        RECT  2.320 1.930 2.930 2.050 ;
        RECT  2.930 1.930 2.960 2.100 ;
        RECT  2.960 1.370 3.120 2.100 ;
        RECT  3.120 1.930 3.150 2.100 ;
        RECT  3.150 1.930 3.760 2.050 ;
        RECT  3.760 1.930 3.790 2.100 ;
        RECT  3.790 1.390 3.950 2.100 ;
        RECT  3.950 1.960 3.980 2.100 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.910 0.725 4.070 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.560 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.155 0.300 ;
        RECT  0.155 -0.300 0.375 0.340 ;
        RECT  0.375 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.860 2.820 ;
        RECT  0.860 2.180 1.080 2.820 ;
        RECT  1.080 2.220 1.680 2.820 ;
        RECT  1.680 2.180 1.900 2.820 ;
        RECT  1.900 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 3.340 2.820 ;
        RECT  3.340 2.180 3.560 2.820 ;
        RECT  3.560 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.800 1.080 1.240 1.240 ;
        RECT  0.680 0.420 0.800 1.660 ;
        RECT  0.550 0.420 0.680 0.580 ;
        RECT  2.470 0.420 2.690 0.590 ;
        RECT  1.930 0.470 2.470 0.590 ;
        RECT  1.710 0.470 1.930 0.885 ;
        RECT  1.150 0.470 1.710 0.590 ;
        RECT  3.170 0.710 3.360 0.870 ;
        RECT  3.050 0.710 3.170 1.190 ;
        RECT  2.620 1.070 3.050 1.190 ;
        RECT  2.500 0.710 2.620 1.190 ;
        RECT  4.190 0.470 4.410 0.890 ;
        RECT  3.720 0.470 4.190 0.590 ;
        RECT  3.500 0.470 3.720 0.885 ;
        RECT  2.930 0.470 3.500 0.590 ;
        RECT  2.810 0.470 2.930 0.950 ;
        RECT  2.070 0.710 2.500 0.870 ;
        RECT  2.770 0.730 2.810 0.950 ;
        RECT  0.930 0.470 1.150 0.890 ;
        RECT  0.420 1.500 0.680 1.660 ;
    END
END IND4D2

MACRO IND4D4
    CLASS CORE ;
    FOREIGN IND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.610 6.030 1.990 ;
        RECT  6.030 0.760 6.450 1.990 ;
        RECT  6.450 1.610 7.160 1.990 ;
        RECT  6.450 0.760 7.260 0.920 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 1.005 7.590 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.900 2.820 ;
        RECT  0.900 2.180 1.120 2.820 ;
        RECT  1.120 2.220 1.700 2.820 ;
        RECT  1.700 2.180 1.920 2.820 ;
        RECT  1.920 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 3.325 2.820 ;
        RECT  3.325 2.180 3.545 2.820 ;
        RECT  3.545 2.220 4.130 2.820 ;
        RECT  4.130 2.180 4.350 2.820 ;
        RECT  4.350 2.220 4.940 2.820 ;
        RECT  4.940 2.180 5.160 2.820 ;
        RECT  5.160 2.220 5.750 2.820 ;
        RECT  5.750 2.180 5.970 2.820 ;
        RECT  5.970 2.220 6.540 2.820 ;
        RECT  6.540 2.180 6.760 2.820 ;
        RECT  6.760 2.220 7.330 2.820 ;
        RECT  7.330 2.180 7.550 2.820 ;
        RECT  7.550 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.700 1.080 2.100 1.240 ;
        RECT  0.700 1.960 0.730 2.100 ;
        RECT  0.610 1.080 0.700 2.100 ;
        RECT  0.540 0.420 0.610 2.100 ;
        RECT  0.450 0.420 0.540 1.240 ;
        RECT  2.720 0.470 4.240 0.630 ;
        RECT  2.500 0.470 2.720 0.890 ;
        RECT  2.000 0.470 2.500 0.590 ;
        RECT  1.780 0.470 2.000 0.890 ;
        RECT  1.280 0.470 1.780 0.590 ;
        RECT  7.400 0.470 7.620 0.885 ;
        RECT  4.360 0.470 7.400 0.630 ;
        RECT  2.860 0.750 5.740 0.885 ;
        RECT  1.060 0.470 1.280 0.890 ;
        RECT  0.510 1.960 0.540 2.100 ;
        LAYER M1 ;
        RECT  1.290 1.610 5.815 1.990 ;
        RECT  6.665 0.760 7.260 0.920 ;
        RECT  6.665 1.610 7.160 1.990 ;
    END
END IND4D4

MACRO INR2D0
    CLASS CORE ;
    FOREIGN INR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.900 1.370 2.060 ;
        RECT  0.840 0.470 1.370 0.630 ;
        RECT  1.370 0.470 1.510 2.060 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.900 1.240 ;
        RECT  0.420 0.470 0.540 2.060 ;
        RECT  0.060 0.470 0.420 0.630 ;
        RECT  0.060 1.900 0.420 2.060 ;
    END
END INR2D0

MACRO INR2D1
    CLASS CORE ;
    FOREIGN INR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.860 0.430 1.080 0.845 ;
        RECT  1.150 1.640 1.370 2.060 ;
        RECT  1.080 0.725 1.370 0.845 ;
        RECT  1.370 0.725 1.510 1.760 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.580 0.710 0.700 1.810 ;
        RECT  0.700 1.080 0.910 1.240 ;
        RECT  0.070 0.710 0.580 0.870 ;
        RECT  0.070 1.650 0.580 1.810 ;
    END
END INR2D1

MACRO INR2D2
    CLASS CORE ;
    FOREIGN INR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.470 1.030 0.885 ;
        RECT  1.130 1.640 1.370 1.800 ;
        RECT  1.030 0.765 1.370 0.885 ;
        RECT  1.370 0.765 1.510 1.800 ;
        RECT  1.510 0.765 1.540 0.890 ;
        RECT  1.540 0.470 1.760 0.890 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 1.810 2.820 ;
        RECT  1.810 2.180 2.030 2.820 ;
        RECT  2.030 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.680 1.030 1.840 2.050 ;
        RECT  0.540 1.930 1.680 2.050 ;
        RECT  0.540 1.080 0.900 1.240 ;
        RECT  0.420 0.710 0.540 2.050 ;
        RECT  0.290 0.710 0.420 0.870 ;
        RECT  0.070 1.640 0.420 2.050 ;
        RECT  0.070 0.470 0.290 0.870 ;
    END
END INR2D2

MACRO INR2D4
    CLASS CORE ;
    FOREIGN INR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.630 1.760 2.050 ;
        RECT  1.760 1.890 3.150 2.050 ;
        RECT  3.150 1.425 3.570 2.050 ;
        RECT  3.570 1.425 3.650 1.565 ;
        RECT  1.090 0.470 3.650 0.630 ;
        RECT  3.650 0.470 3.770 1.565 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.710 1.235 ;
        RECT  1.710 1.005 1.830 1.510 ;
        RECT  1.830 1.390 2.770 1.510 ;
        RECT  2.770 1.030 2.930 1.510 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 3.490 2.820 ;
        RECT  3.490 2.180 3.710 2.820 ;
        RECT  3.710 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.360 0.750 3.520 1.255 ;
        RECT  2.390 0.750 3.360 0.885 ;
        RECT  2.230 0.750 2.390 1.270 ;
        RECT  1.200 0.750 2.230 0.885 ;
        RECT  1.080 0.750 1.200 1.240 ;
        RECT  0.670 1.080 1.080 1.240 ;
        RECT  0.670 1.960 0.700 2.100 ;
        RECT  0.610 1.080 0.670 2.100 ;
        RECT  0.510 0.420 0.610 2.100 ;
        RECT  0.450 0.420 0.510 1.240 ;
        RECT  0.480 1.960 0.510 2.100 ;
        LAYER M1 ;
        RECT  3.650 0.470 3.770 1.210 ;
        RECT  1.760 1.890 2.935 2.050 ;
        RECT  1.540 1.630 1.760 2.050 ;
        RECT  1.090 0.470 3.650 0.630 ;
    END
END INR2D4

MACRO INR3D0
    CLASS CORE ;
    FOREIGN INR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.810 0.470 1.660 0.630 ;
        RECT  1.480 1.635 1.690 2.050 ;
        RECT  1.660 0.470 1.690 0.690 ;
        RECT  1.690 0.470 1.700 2.050 ;
        RECT  1.700 0.470 1.830 1.755 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.230 0.300 ;
        RECT  1.230 -0.300 1.450 0.340 ;
        RECT  1.450 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.090 0.910 1.250 ;
        RECT  0.420 0.480 0.540 1.800 ;
        RECT  0.070 0.480 0.420 0.640 ;
        RECT  0.070 1.640 0.420 1.800 ;
    END
END INR3D0

MACRO INR3D1
    CLASS CORE ;
    FOREIGN INR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.750 0.710 1.370 0.870 ;
        RECT  1.370 0.710 1.510 1.800 ;
        RECT  1.510 1.640 1.700 1.800 ;
        RECT  1.510 0.710 1.750 0.870 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.030 1.170 2.040 ;
        RECT  1.170 1.920 2.010 2.040 ;
        RECT  1.870 0.730 2.010 0.885 ;
        RECT  2.010 0.730 2.150 2.040 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.140 0.300 ;
        RECT  1.140 -0.300 1.360 0.340 ;
        RECT  1.360 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 2.400 2.820 ;
        RECT  2.400 2.180 2.620 2.820 ;
        RECT  2.620 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.230 0.430 2.470 0.590 ;
        RECT  0.630 0.470 2.230 0.590 ;
        RECT  0.630 1.080 0.870 1.240 ;
        RECT  0.510 0.470 0.630 1.780 ;
        RECT  0.280 0.765 0.510 0.885 ;
        RECT  0.280 1.640 0.510 1.780 ;
        RECT  0.060 0.470 0.280 0.885 ;
        RECT  0.060 1.640 0.280 2.060 ;
    END
END INR3D1

MACRO INR3D2
    CLASS CORE ;
    FOREIGN INR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 0.470 1.010 0.900 ;
        RECT  1.010 0.470 1.510 0.590 ;
        RECT  1.510 0.470 1.730 0.885 ;
        RECT  1.730 0.470 2.220 0.590 ;
        RECT  2.220 0.470 2.440 0.900 ;
        RECT  1.530 1.890 2.650 2.050 ;
        RECT  2.440 0.780 2.650 0.900 ;
        RECT  2.650 0.780 2.790 2.050 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.030 1.180 1.515 ;
        RECT  1.180 1.395 2.010 1.515 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.080 2.250 1.240 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 2.520 2.820 ;
        RECT  2.520 2.180 2.740 2.820 ;
        RECT  2.740 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.070 0.470 0.290 0.870 ;
        RECT  0.290 1.640 0.435 1.770 ;
        RECT  0.290 0.710 0.435 0.870 ;
        RECT  0.435 0.710 0.555 1.770 ;
        RECT  0.555 1.080 0.890 1.240 ;
        RECT  0.555 1.650 2.380 1.770 ;
        RECT  2.380 1.050 2.530 1.770 ;
        RECT  0.070 1.640 0.290 2.040 ;
    END
END INR3D2

MACRO INR3D4
    CLASS CORE ;
    FOREIGN INR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.430 1.330 0.590 ;
        RECT  1.330 0.470 1.800 0.590 ;
        RECT  1.800 0.430 2.020 0.590 ;
        RECT  2.020 0.470 2.490 0.590 ;
        RECT  2.490 0.430 2.710 0.590 ;
        RECT  2.710 0.470 3.180 0.590 ;
        RECT  3.180 0.430 3.400 0.590 ;
        RECT  1.780 1.890 3.870 2.050 ;
        RECT  3.400 0.470 3.870 0.590 ;
        RECT  3.870 1.650 4.090 2.050 ;
        RECT  3.870 0.430 4.090 0.590 ;
        RECT  4.090 1.890 4.430 2.050 ;
        RECT  4.090 0.470 4.560 0.590 ;
        RECT  4.560 0.430 4.780 0.590 ;
        RECT  4.430 1.425 4.850 2.050 ;
        RECT  4.850 1.425 4.990 1.545 ;
        RECT  4.780 0.470 4.990 0.590 ;
        RECT  4.990 0.470 5.110 1.545 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.950 1.840 1.515 ;
        RECT  1.840 0.950 2.610 1.070 ;
        RECT  2.610 0.950 2.730 1.515 ;
        RECT  2.730 1.395 3.130 1.515 ;
        RECT  3.130 0.950 3.250 1.515 ;
        RECT  3.250 0.950 3.790 1.070 ;
        RECT  3.790 0.950 3.950 1.285 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.095 1.370 1.255 ;
        RECT  1.370 1.005 1.520 1.755 ;
        RECT  1.520 1.635 2.270 1.755 ;
        RECT  2.270 1.190 2.490 1.755 ;
        RECT  2.490 1.635 3.370 1.755 ;
        RECT  3.370 1.190 3.590 1.755 ;
        RECT  3.590 1.410 4.095 1.530 ;
        RECT  4.095 1.035 4.215 1.530 ;
        RECT  4.215 1.035 4.235 1.255 ;
        RECT  4.235 1.035 4.580 1.195 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.970 0.300 ;
        RECT  4.970 -0.300 5.190 0.340 ;
        RECT  5.190 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.780 2.820 ;
        RECT  2.780 2.180 3.000 2.820 ;
        RECT  3.000 2.220 4.830 2.820 ;
        RECT  4.830 2.180 5.050 2.820 ;
        RECT  5.050 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.020 0.710 1.180 1.800 ;
        RECT  1.180 0.710 2.850 0.830 ;
        RECT  2.850 0.710 3.010 1.275 ;
        RECT  3.010 0.710 4.710 0.830 ;
        RECT  4.710 0.710 4.870 1.245 ;
        RECT  0.640 0.710 1.020 0.870 ;
        RECT  0.710 1.640 1.020 1.800 ;
        RECT  0.490 1.640 0.710 2.060 ;
        RECT  0.420 0.450 0.640 0.870 ;
        LAYER M1 ;
        RECT  1.090 0.430 1.330 0.590 ;
        RECT  1.780 1.890 3.870 2.050 ;
        RECT  3.870 1.650 4.090 2.050 ;
        RECT  4.090 1.890 4.215 2.050 ;
        RECT  1.330 0.470 1.800 0.590 ;
        RECT  1.800 0.430 2.020 0.590 ;
        RECT  2.020 0.470 2.490 0.590 ;
        RECT  2.490 0.430 2.710 0.590 ;
        RECT  2.710 0.470 3.180 0.590 ;
        RECT  3.180 0.430 3.400 0.590 ;
        RECT  3.400 0.470 3.870 0.590 ;
        RECT  3.870 0.430 4.090 0.590 ;
        RECT  4.090 0.470 4.560 0.590 ;
        RECT  4.560 0.430 4.780 0.590 ;
        RECT  4.780 0.470 4.990 0.590 ;
        RECT  4.990 0.470 5.110 1.210 ;
    END
END INR3D4

MACRO INR4D0
    CLASS CORE ;
    FOREIGN INR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.640 2.010 2.060 ;
        RECT  0.790 0.610 2.010 0.770 ;
        RECT  2.010 0.610 2.050 2.060 ;
        RECT  2.050 0.610 2.150 1.760 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.550 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.180 0.300 ;
        RECT  1.180 -0.300 1.400 0.340 ;
        RECT  1.400 -0.300 1.890 0.300 ;
        RECT  1.890 -0.300 2.110 0.340 ;
        RECT  2.110 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.910 1.240 ;
        RECT  0.420 0.560 0.540 1.800 ;
        RECT  0.070 0.560 0.420 0.720 ;
        RECT  0.070 1.640 0.420 1.800 ;
    END
END INR4D0

MACRO INR4D1
    CLASS CORE ;
    FOREIGN INR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.400 2.820 1.810 ;
        RECT  2.820 1.400 2.970 1.560 ;
        RECT  1.610 0.725 2.970 0.885 ;
        RECT  2.970 0.725 3.110 1.560 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.270 0.725 3.430 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END B3
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.820 ;
        RECT  1.470 -0.300 2.800 0.300 ;
        RECT  2.800 -0.300 3.020 0.605 ;
        RECT  3.020 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.750 1.080 1.560 1.240 ;
        RECT  0.660 0.450 0.750 1.240 ;
        RECT  0.590 0.450 0.660 1.850 ;
        RECT  3.420 1.960 3.450 2.100 ;
        RECT  3.260 1.390 3.420 2.100 ;
        RECT  3.230 1.930 3.260 2.100 ;
        RECT  1.030 1.930 3.230 2.050 ;
        RECT  1.000 1.930 1.030 2.100 ;
        RECT  0.840 1.370 1.000 2.100 ;
        RECT  0.500 1.080 0.590 1.850 ;
        RECT  0.810 1.930 0.840 2.100 ;
    END
END INR4D1

MACRO INR4D2
    CLASS CORE ;
    FOREIGN INR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.900 1.390 6.120 1.810 ;
        RECT  6.120 1.390 6.490 1.510 ;
        RECT  1.740 0.530 6.490 0.690 ;
        RECT  6.490 0.530 6.630 1.510 ;
        RECT  6.630 1.390 6.660 1.510 ;
        RECT  6.660 1.390 6.880 1.810 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.520 0.300 ;
        RECT  0.520 -0.300 0.740 0.340 ;
        RECT  0.740 -0.300 1.350 0.300 ;
        RECT  1.350 -0.300 1.570 0.340 ;
        RECT  1.570 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.340 ;
        RECT  2.390 -0.300 2.870 0.300 ;
        RECT  2.870 -0.300 3.090 0.340 ;
        RECT  3.090 -0.300 3.690 0.300 ;
        RECT  3.690 -0.300 3.910 0.340 ;
        RECT  3.910 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.340 ;
        RECT  4.460 -0.300 5.060 0.300 ;
        RECT  5.060 -0.300 5.280 0.340 ;
        RECT  5.280 -0.300 5.610 0.300 ;
        RECT  5.610 -0.300 5.830 0.340 ;
        RECT  5.830 -0.300 6.430 0.300 ;
        RECT  6.430 -0.300 6.650 0.340 ;
        RECT  6.650 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.610 1.010 1.890 1.170 ;
        RECT  0.610 1.930 0.640 2.090 ;
        RECT  0.450 0.740 0.610 2.090 ;
        RECT  0.330 0.740 0.450 0.860 ;
        RECT  0.420 1.930 0.450 2.090 ;
        RECT  3.850 1.960 3.880 2.100 ;
        RECT  3.690 1.390 3.850 2.100 ;
        RECT  3.660 1.930 3.690 2.100 ;
        RECT  3.120 1.930 3.660 2.050 ;
        RECT  2.900 1.630 3.120 2.050 ;
        RECT  2.360 1.930 2.900 2.050 ;
        RECT  2.330 1.930 2.360 2.100 ;
        RECT  2.170 1.370 2.330 2.100 ;
        RECT  2.140 1.930 2.170 2.100 ;
        RECT  1.670 1.930 2.140 2.050 ;
        RECT  1.640 1.930 1.670 2.100 ;
        RECT  1.480 1.370 1.640 2.100 ;
        RECT  1.450 1.930 1.480 2.100 ;
        RECT  0.980 1.930 1.450 2.050 ;
        RECT  0.950 1.930 0.980 2.100 ;
        RECT  0.790 1.370 0.950 2.100 ;
        RECT  5.140 1.390 5.360 1.810 ;
        RECT  4.600 1.390 5.140 1.510 ;
        RECT  4.500 1.390 4.600 1.810 ;
        RECT  4.380 1.150 4.500 1.810 ;
        RECT  3.500 1.150 4.380 1.270 ;
        RECT  3.380 1.150 3.500 1.810 ;
        RECT  3.280 1.390 3.380 1.810 ;
        RECT  2.740 1.390 3.280 1.510 ;
        RECT  7.230 1.960 7.260 2.100 ;
        RECT  7.070 1.370 7.230 2.100 ;
        RECT  7.040 1.930 7.070 2.100 ;
        RECT  6.500 1.930 7.040 2.050 ;
        RECT  6.280 1.630 6.500 2.050 ;
        RECT  5.740 1.930 6.280 2.050 ;
        RECT  5.710 1.930 5.740 2.100 ;
        RECT  5.550 1.370 5.710 2.100 ;
        RECT  5.520 1.930 5.550 2.100 ;
        RECT  4.980 1.930 5.520 2.050 ;
        RECT  4.760 1.630 4.980 2.050 ;
        RECT  4.220 1.930 4.760 2.050 ;
        RECT  4.190 1.930 4.220 2.100 ;
        RECT  4.030 1.390 4.190 2.100 ;
        RECT  4.000 1.960 4.030 2.100 ;
        RECT  2.520 1.390 2.740 1.810 ;
        RECT  0.760 1.960 0.790 2.100 ;
        RECT  0.110 0.440 0.330 0.860 ;
    END
END INR4D2

MACRO INR4D4
    CLASS CORE ;
    FOREIGN INR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.240 1.560 6.670 1.720 ;
        RECT  1.290 0.490 6.670 0.870 ;
        RECT  6.670 0.490 7.090 1.720 ;
        RECT  7.090 0.490 7.170 0.870 ;
        RECT  7.090 1.560 7.260 1.720 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 0.900 0.300 ;
        RECT  0.900 -0.300 1.120 0.340 ;
        RECT  1.120 -0.300 1.690 0.300 ;
        RECT  1.690 -0.300 1.910 0.340 ;
        RECT  1.910 -0.300 2.500 0.300 ;
        RECT  2.500 -0.300 2.720 0.340 ;
        RECT  2.720 -0.300 3.310 0.300 ;
        RECT  3.310 -0.300 3.530 0.340 ;
        RECT  3.530 -0.300 4.130 0.300 ;
        RECT  4.130 -0.300 4.350 0.340 ;
        RECT  4.350 -0.300 4.950 0.300 ;
        RECT  4.950 -0.300 5.170 0.340 ;
        RECT  5.170 -0.300 5.760 0.300 ;
        RECT  5.760 -0.300 5.980 0.340 ;
        RECT  5.980 -0.300 6.560 0.300 ;
        RECT  6.560 -0.300 6.780 0.340 ;
        RECT  6.780 -0.300 7.340 0.300 ;
        RECT  7.340 -0.300 7.560 0.340 ;
        RECT  7.560 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.700 1.080 2.230 1.240 ;
        RECT  0.610 0.420 0.700 1.240 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.540 0.420 0.610 2.100 ;
        RECT  0.450 1.080 0.540 2.100 ;
        RECT  2.720 1.890 4.240 2.050 ;
        RECT  2.690 1.890 2.720 2.100 ;
        RECT  2.530 1.370 2.690 2.100 ;
        RECT  2.500 1.930 2.530 2.100 ;
        RECT  2.000 1.930 2.500 2.050 ;
        RECT  1.970 1.930 2.000 2.100 ;
        RECT  1.810 1.370 1.970 2.100 ;
        RECT  1.780 1.930 1.810 2.100 ;
        RECT  1.280 1.930 1.780 2.050 ;
        RECT  1.250 1.930 1.280 2.100 ;
        RECT  1.090 1.370 1.250 2.100 ;
        RECT  7.430 1.550 7.590 2.050 ;
        RECT  6.100 1.890 7.430 2.050 ;
        RECT  6.070 1.890 6.100 2.100 ;
        RECT  5.910 1.370 6.070 2.100 ;
        RECT  5.880 1.890 5.910 2.100 ;
        RECT  4.360 1.890 5.880 2.050 ;
        RECT  2.860 1.610 5.740 1.770 ;
        RECT  1.060 1.960 1.090 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
        LAYER M1 ;
        RECT  1.290 0.490 6.455 0.870 ;
        RECT  6.240 1.560 6.455 1.720 ;
    END
END INR4D4

MACRO INVD0
    CLASS CORE ;
    FOREIGN INVD0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.660 0.550 1.710 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.640 2.820 ;
        END
    END VDD
END INVD0

MACRO INVD1
    CLASS CORE ;
    FOREIGN INVD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.960 0.390 2.100 ;
        RECT  0.390 0.420 0.550 2.100 ;
        RECT  0.550 1.960 0.580 2.100 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
END INVD1

MACRO INVD12
    CLASS CORE ;
    FOREIGN INVD12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.640 2.190 2.020 ;
        RECT  0.460 0.500 2.190 0.880 ;
        RECT  2.190 0.500 2.610 2.020 ;
        RECT  2.610 1.640 4.330 2.020 ;
        RECT  2.610 0.500 4.330 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        RECT  0.230 1.080 1.030 1.240 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.460 0.500 1.975 0.880 ;
        RECT  0.460 1.640 1.975 2.020 ;
        RECT  2.825 0.500 4.330 0.880 ;
        RECT  2.825 1.640 4.330 2.020 ;
    END
END INVD12

MACRO INVD16
    CLASS CORE ;
    FOREIGN INVD16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 2.830 2.020 ;
        RECT  0.440 0.500 2.830 0.880 ;
        RECT  2.830 0.500 3.250 2.020 ;
        RECT  3.250 1.640 5.640 2.020 ;
        RECT  3.250 0.500 5.640 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        RECT  0.230 1.080 0.980 1.240 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.440 0.500 2.615 0.880 ;
        RECT  0.440 1.640 2.615 2.020 ;
        RECT  3.465 0.500 5.640 0.880 ;
        RECT  3.465 1.640 5.640 2.020 ;
    END
END INVD16

MACRO INVD2
    CLASS CORE ;
    FOREIGN INVD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.960 0.400 2.100 ;
        RECT  0.400 0.420 0.560 2.100 ;
        RECT  0.560 1.960 0.590 2.100 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.960 2.820 ;
        END
    END VDD
END INVD2

MACRO INVD20
    CLASS CORE ;
    FOREIGN INVD20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.640 3.470 2.020 ;
        RECT  0.420 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 6.940 2.020 ;
        RECT  3.890 0.500 6.940 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        RECT  0.230 1.080 0.990 1.240 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.420 0.500 3.255 0.880 ;
        RECT  0.420 1.640 3.255 2.020 ;
        RECT  4.105 0.500 6.940 0.880 ;
        RECT  4.105 1.640 6.940 2.020 ;
    END
END INVD20

MACRO INVD24
    CLASS CORE ;
    FOREIGN INVD24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 4.110 2.020 ;
        RECT  0.440 0.500 4.110 0.880 ;
        RECT  4.110 0.500 4.530 2.020 ;
        RECT  4.530 1.640 8.520 2.020 ;
        RECT  4.530 0.500 8.520 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.080 1.000 1.240 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.440 0.500 3.895 0.880 ;
        RECT  0.440 1.640 3.895 2.020 ;
        RECT  4.745 0.500 8.520 0.880 ;
        RECT  4.745 1.640 8.520 2.020 ;
    END
END INVD24

MACRO INVD3
    CLASS CORE ;
    FOREIGN INVD3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.640 0.590 2.020 ;
        RECT  0.520 0.500 0.590 0.880 ;
        RECT  0.590 0.500 1.010 2.020 ;
        RECT  1.010 1.640 1.530 2.020 ;
        RECT  1.010 0.500 1.530 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.910 0.300 ;
        RECT  0.910 -0.300 1.130 0.340 ;
        RECT  1.130 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.910 2.820 ;
        RECT  0.910 2.180 1.130 2.820 ;
        RECT  1.130 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.225 0.500 1.530 0.880 ;
        RECT  1.225 1.640 1.530 2.020 ;
    END
END INVD3

MACRO INVD4
    CLASS CORE ;
    FOREIGN INVD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.640 0.910 2.020 ;
        RECT  0.470 0.500 0.910 0.880 ;
        RECT  0.910 0.500 1.330 2.020 ;
        RECT  1.330 1.640 1.440 2.020 ;
        RECT  1.330 0.500 1.440 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.470 0.500 0.695 0.880 ;
        RECT  0.470 1.640 0.695 2.020 ;
    END
END INVD4

MACRO INVD6
    CLASS CORE ;
    FOREIGN INVD6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.640 0.910 2.020 ;
        RECT  0.450 0.500 0.910 0.880 ;
        RECT  0.910 0.500 1.330 2.020 ;
        RECT  1.330 1.640 2.110 2.020 ;
        RECT  1.330 0.500 2.110 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.450 0.500 0.695 0.880 ;
        RECT  0.450 1.640 0.695 2.020 ;
        RECT  1.545 0.500 2.110 0.880 ;
        RECT  1.545 1.640 2.110 2.020 ;
    END
END INVD6

MACRO INVD8
    CLASS CORE ;
    FOREIGN INVD8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.640 1.230 2.020 ;
        RECT  0.440 0.500 1.230 0.880 ;
        RECT  1.230 0.500 1.650 2.020 ;
        RECT  1.650 1.640 2.770 2.020 ;
        RECT  1.650 0.500 2.770 0.880 ;
        END
    END ZN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.440 0.500 1.015 0.880 ;
        RECT  0.440 1.640 1.015 2.020 ;
        RECT  1.865 0.500 2.770 0.880 ;
        RECT  1.865 1.640 2.770 2.020 ;
    END
END INVD8

MACRO IOA21D0
    CLASS CORE ;
    FOREIGN IOA21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.890 1.690 2.050 ;
        RECT  1.470 0.470 1.690 0.630 ;
        RECT  1.690 0.470 1.830 2.050 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.830 0.300 ;
        RECT  0.830 -0.300 1.050 0.340 ;
        RECT  1.050 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.520 1.200 1.770 ;
        RECT  0.140 0.520 1.040 0.680 ;
        RECT  0.660 1.650 1.040 1.770 ;
        RECT  0.500 1.650 0.660 2.010 ;
    END
END IOA21D0

MACRO IOA21D1
    CLASS CORE ;
    FOREIGN IOA21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.890 1.690 2.050 ;
        RECT  1.490 0.420 1.690 0.840 ;
        RECT  1.690 0.420 1.710 2.050 ;
        RECT  1.710 0.720 1.830 2.050 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.830 0.300 ;
        RECT  0.830 -0.300 1.050 0.340 ;
        RECT  1.050 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.040 0.470 1.200 1.770 ;
        RECT  0.140 0.470 1.040 0.630 ;
        RECT  0.660 1.650 1.040 1.770 ;
        RECT  0.500 1.650 0.660 2.090 ;
    END
END IOA21D1

MACRO IOA21D2
    CLASS CORE ;
    FOREIGN IOA21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.200 1.960 1.230 2.100 ;
        RECT  1.230 1.390 1.390 2.100 ;
        RECT  1.390 1.960 1.420 2.100 ;
        RECT  1.390 0.710 1.510 1.510 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.950 1.390 2.010 2.100 ;
        RECT  1.510 0.710 2.010 0.870 ;
        RECT  2.010 0.710 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.710 2.150 1.515 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.810 2.820 ;
        RECT  0.810 2.180 1.030 2.820 ;
        RECT  1.030 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.470 2.430 1.290 ;
        RECT  1.260 0.470 2.270 0.590 ;
        RECT  1.100 0.470 1.260 1.270 ;
        RECT  0.890 0.470 1.100 0.590 ;
        RECT  0.670 0.470 0.890 0.885 ;
        RECT  0.610 0.765 0.670 0.885 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.450 0.765 0.610 2.100 ;
        RECT  0.420 1.960 0.450 2.100 ;
    END
END IOA21D2

MACRO IOA21D4
    CLASS CORE ;
    FOREIGN IOA21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.650 1.230 2.030 ;
        RECT  1.230 1.425 1.380 2.030 ;
        RECT  1.380 0.710 1.500 2.030 ;
        RECT  1.500 1.425 1.650 2.030 ;
        RECT  1.500 0.710 1.720 0.870 ;
        RECT  1.650 1.650 3.030 2.030 ;
        RECT  2.830 0.710 3.030 0.870 ;
        RECT  3.030 0.710 3.150 2.030 ;
        RECT  3.150 1.650 3.410 2.030 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.140 1.080 2.260 1.240 ;
        RECT  2.260 0.470 2.380 1.240 ;
        RECT  2.380 0.470 3.290 0.590 ;
        RECT  3.290 0.470 3.430 1.235 ;
        RECT  3.430 1.075 3.570 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.080 0.730 1.240 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.750 0.300 ;
        RECT  0.750 -0.300 0.970 0.340 ;
        RECT  0.970 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 3.490 0.300 ;
        RECT  3.490 -0.300 3.710 0.340 ;
        RECT  3.710 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.750 1.030 2.910 1.480 ;
        RECT  1.990 1.360 2.750 1.480 ;
        RECT  1.870 0.470 1.990 1.480 ;
        RECT  0.870 0.470 1.870 0.590 ;
        RECT  1.630 1.040 1.870 1.200 ;
        RECT  0.750 0.470 0.870 0.885 ;
        RECT  0.490 0.765 0.750 0.885 ;
        RECT  0.610 1.960 0.640 2.100 ;
        RECT  0.490 1.390 0.610 2.100 ;
        RECT  0.450 0.765 0.490 2.100 ;
        RECT  0.370 0.765 0.450 1.510 ;
        RECT  0.420 1.960 0.450 2.100 ;
        RECT  0.310 0.765 0.370 0.885 ;
        RECT  0.090 0.470 0.310 0.885 ;
        LAYER M1 ;
        RECT  1.865 1.650 3.030 2.030 ;
        RECT  1.380 0.710 1.500 1.210 ;
        RECT  1.500 0.710 1.720 0.870 ;
        RECT  2.830 0.710 3.030 0.870 ;
        RECT  3.030 0.710 3.150 2.030 ;
        RECT  3.150 1.650 3.410 2.030 ;
    END
END IOA21D4

MACRO IOA22D0
    CLASS CORE ;
    FOREIGN IOA22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.890 1.050 2.050 ;
        RECT  0.950 0.710 1.050 0.870 ;
        RECT  1.050 0.710 1.190 2.050 ;
        RECT  1.190 1.890 2.170 2.050 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.535 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.535 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.660 0.300 ;
        RECT  1.660 -0.300 1.880 0.870 ;
        RECT  1.880 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.170 0.350 2.820 ;
        RECT  0.350 2.220 0.650 2.820 ;
        RECT  0.650 2.170 0.870 2.820 ;
        RECT  0.870 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 1.090 0.930 1.250 ;
        RECT  0.710 0.660 0.830 1.860 ;
        RECT  0.590 0.660 0.710 0.820 ;
        RECT  0.340 1.700 0.710 1.860 ;
    END
END IOA22D0

MACRO IOA22D1
    CLASS CORE ;
    FOREIGN IOA22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 0.420 1.220 0.900 ;
        RECT  1.240 1.960 1.270 2.100 ;
        RECT  1.220 0.420 1.290 1.125 ;
        RECT  1.290 0.780 1.340 1.125 ;
        RECT  1.270 1.390 1.370 2.100 ;
        RECT  1.340 1.005 1.370 1.125 ;
        RECT  1.370 1.005 1.430 2.100 ;
        RECT  1.430 1.930 1.460 2.100 ;
        RECT  1.430 1.005 1.510 1.515 ;
        RECT  1.460 1.930 2.270 2.050 ;
        RECT  2.270 1.635 2.490 2.050 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.180 0.770 1.400 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 1.870 0.300 ;
        RECT  1.870 -0.300 2.090 0.340 ;
        RECT  2.090 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.900 2.820 ;
        RECT  0.900 2.180 1.120 2.820 ;
        RECT  1.120 2.220 1.630 2.820 ;
        RECT  1.630 2.180 1.850 2.820 ;
        RECT  1.850 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.010 1.050 1.100 1.270 ;
        RECT  0.890 0.650 1.010 2.050 ;
        RECT  0.740 0.650 0.890 0.810 ;
        RECT  2.270 0.470 2.490 0.885 ;
        RECT  1.700 0.470 2.270 0.590 ;
        RECT  0.490 1.890 0.890 2.050 ;
        RECT  1.480 0.470 1.700 0.885 ;
    END
END IOA22D1

MACRO IOA22D2
    CLASS CORE ;
    FOREIGN IOA22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.910 1.960 1.940 2.100 ;
        RECT  1.940 1.390 2.010 2.100 ;
        RECT  1.620 0.710 2.010 0.870 ;
        RECT  2.010 0.710 2.100 2.100 ;
        RECT  2.100 1.960 2.130 2.100 ;
        RECT  2.100 0.710 2.150 1.515 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.060 2.590 1.280 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 0.725 3.110 1.255 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 1.210 0.300 ;
        RECT  1.210 -0.300 1.430 0.340 ;
        RECT  1.430 -0.300 2.030 0.300 ;
        RECT  2.030 -0.300 2.250 0.340 ;
        RECT  2.250 -0.300 2.850 0.300 ;
        RECT  2.850 -0.300 3.070 0.340 ;
        RECT  3.070 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.260 1.390 0.480 1.510 ;
        RECT  0.480 0.710 0.600 1.510 ;
        RECT  0.600 0.710 1.380 0.870 ;
        RECT  1.380 0.710 1.500 1.240 ;
        RECT  1.500 1.080 1.850 1.240 ;
        RECT  0.670 1.660 1.200 1.780 ;
        RECT  1.200 1.660 1.420 2.090 ;
        RECT  0.100 1.390 0.260 2.100 ;
        RECT  3.100 1.960 3.130 2.100 ;
        RECT  2.940 1.390 3.100 2.100 ;
        RECT  2.830 1.390 2.940 1.510 ;
        RECT  2.910 1.960 2.940 2.100 ;
        RECT  2.710 0.470 2.830 1.510 ;
        RECT  2.450 0.470 2.710 0.630 ;
        RECT  0.360 0.470 2.450 0.590 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.200 0.470 0.360 1.270 ;
        RECT  0.450 1.660 0.670 2.090 ;
    END
END IOA22D2

MACRO IOA22D4
    CLASS CORE ;
    FOREIGN IOA22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.625 1.650 3.790 2.030 ;
        RECT  3.625 0.490 3.790 0.870 ;
        RECT  3.790 0.490 4.210 2.030 ;
        RECT  4.210 0.490 4.590 0.870 ;
        RECT  4.210 1.650 4.600 2.030 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.110 1.515 ;
        RECT  3.110 1.050 3.245 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.640 1.005 2.800 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        RECT  0.240 1.395 1.265 1.515 ;
        RECT  1.265 1.030 1.425 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.580 0.300 ;
        RECT  2.580 -0.300 2.800 0.340 ;
        RECT  2.800 -0.300 3.225 0.300 ;
        RECT  3.225 -0.300 3.445 0.340 ;
        RECT  3.445 -0.300 4.770 0.300 ;
        RECT  4.770 -0.300 4.990 0.340 ;
        RECT  4.990 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.225 2.820 ;
        RECT  3.225 2.180 3.445 2.820 ;
        RECT  3.445 2.220 4.770 2.820 ;
        RECT  4.770 2.180 4.990 2.820 ;
        RECT  4.990 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.985 1.930 2.455 2.050 ;
        RECT  0.765 1.670 0.985 2.050 ;
        RECT  0.290 1.930 0.765 2.050 ;
        RECT  2.325 0.720 3.110 0.880 ;
        RECT  2.575 1.650 2.795 2.050 ;
        RECT  2.325 1.650 2.575 1.810 ;
        RECT  2.205 0.720 2.325 1.810 ;
        RECT  3.505 1.050 3.570 1.270 ;
        RECT  3.385 0.470 3.505 1.270 ;
        RECT  1.710 0.470 3.385 0.590 ;
        RECT  1.710 1.650 2.075 1.810 ;
        RECT  1.550 0.470 1.710 1.810 ;
        RECT  0.290 0.470 1.550 0.590 ;
        RECT  1.880 1.080 2.205 1.240 ;
        RECT  0.070 1.670 0.290 2.050 ;
        RECT  0.070 0.470 0.290 0.870 ;
        RECT  0.430 0.710 1.380 0.870 ;
        LAYER M1 ;
        RECT  4.425 0.490 4.590 0.870 ;
        RECT  4.425 1.650 4.600 2.030 ;
    END
END IOA22D4

MACRO LHCND1
    CLASS CORE ;
    FOREIGN LHCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.940 3.830 2.100 ;
        RECT  3.830 1.390 3.930 2.100 ;
        RECT  3.780 0.710 3.930 0.870 ;
        RECT  3.930 0.710 3.990 2.100 ;
        RECT  3.990 1.940 4.020 2.100 ;
        RECT  3.990 0.710 4.070 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.940 4.550 2.100 ;
        RECT  4.550 1.390 4.570 2.100 ;
        RECT  4.550 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.710 2.100 ;
        RECT  4.710 1.940 4.740 2.100 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.395 1.370 1.515 ;
        RECT  1.370 0.880 1.530 1.515 ;
        RECT  1.530 1.355 2.180 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.250 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.250 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 2.370 0.300 ;
        RECT  2.370 -0.300 2.590 0.340 ;
        RECT  2.590 -0.300 3.130 0.300 ;
        RECT  3.130 -0.300 3.350 0.340 ;
        RECT  3.350 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.130 2.820 ;
        RECT  3.130 2.180 3.350 2.820 ;
        RECT  3.350 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 1.930 1.820 2.090 ;
        RECT  0.260 1.930 1.580 2.050 ;
        RECT  2.450 1.080 2.750 1.240 ;
        RECT  2.330 0.580 2.450 1.810 ;
        RECT  1.450 0.580 2.330 0.740 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  2.990 1.050 3.360 1.270 ;
        RECT  2.870 0.480 2.990 2.050 ;
        RECT  2.750 0.480 2.870 0.640 ;
        RECT  2.770 1.630 2.870 2.050 ;
        RECT  2.400 1.930 2.770 2.050 ;
        RECT  4.420 1.050 4.450 1.290 ;
        RECT  4.300 0.470 4.420 1.290 ;
        RECT  3.640 0.470 4.300 0.590 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.050 ;
        RECT  3.480 0.470 3.640 1.830 ;
    END
END LHCND1

MACRO LHCND2
    CLASS CORE ;
    FOREIGN LHCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.790 1.940 3.820 2.100 ;
        RECT  3.820 1.390 3.930 2.100 ;
        RECT  3.770 0.710 3.930 0.870 ;
        RECT  3.930 0.710 3.980 2.100 ;
        RECT  3.980 1.940 4.010 2.100 ;
        RECT  3.980 0.710 4.070 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.940 4.510 2.100 ;
        RECT  4.510 1.390 4.570 2.100 ;
        RECT  4.510 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.670 2.100 ;
        RECT  4.670 1.940 4.700 2.100 ;
        RECT  4.670 0.780 4.710 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.395 1.370 1.515 ;
        RECT  1.370 0.880 1.530 1.515 ;
        RECT  1.530 1.355 2.180 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.250 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.250 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 3.390 0.300 ;
        RECT  3.390 -0.300 3.610 0.340 ;
        RECT  3.610 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.390 2.820 ;
        RECT  3.390 2.180 3.610 2.820 ;
        RECT  3.610 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 1.930 1.820 2.090 ;
        RECT  0.260 1.930 1.580 2.050 ;
        RECT  2.450 1.080 2.720 1.240 ;
        RECT  2.330 0.580 2.450 1.810 ;
        RECT  1.450 0.580 2.330 0.740 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  3.470 1.030 3.630 2.050 ;
        RECT  2.960 1.930 3.470 2.050 ;
        RECT  2.840 0.470 2.960 2.050 ;
        RECT  2.720 0.470 2.840 0.630 ;
        RECT  2.740 1.630 2.840 2.050 ;
        RECT  2.400 1.930 2.740 2.050 ;
        RECT  4.360 1.050 4.430 1.270 ;
        RECT  4.220 0.470 4.360 1.270 ;
        RECT  3.280 0.470 4.220 0.590 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  3.120 0.470 3.280 1.710 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.050 ;
    END
END LHCND2

MACRO LHCND4
    CLASS CORE ;
    FOREIGN LHCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.650 4.110 2.030 ;
        RECT  3.830 0.760 4.110 0.920 ;
        RECT  4.110 0.760 4.530 2.030 ;
        RECT  4.530 1.650 4.800 2.030 ;
        RECT  4.530 0.760 4.820 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.650 5.710 2.030 ;
        RECT  5.310 0.490 5.710 0.870 ;
        RECT  5.710 0.490 6.130 2.030 ;
        RECT  6.130 1.650 6.260 2.030 ;
        RECT  6.130 0.490 6.260 0.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.395 1.370 1.515 ;
        RECT  1.370 0.880 1.530 1.515 ;
        RECT  1.530 1.355 2.180 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.250 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.250 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 3.450 0.300 ;
        RECT  3.450 -0.300 3.670 0.340 ;
        RECT  3.670 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.450 2.820 ;
        RECT  3.450 2.180 3.670 2.820 ;
        RECT  3.670 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 1.930 1.820 2.090 ;
        RECT  0.260 1.930 1.580 2.050 ;
        RECT  2.450 1.080 2.720 1.240 ;
        RECT  2.330 0.580 2.450 1.810 ;
        RECT  1.450 0.580 2.330 0.740 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  3.455 1.030 3.615 2.050 ;
        RECT  2.960 1.930 3.455 2.050 ;
        RECT  2.840 0.470 2.960 2.050 ;
        RECT  2.720 0.470 2.840 0.630 ;
        RECT  2.740 1.630 2.840 2.050 ;
        RECT  2.400 1.930 2.740 2.050 ;
        RECT  5.140 1.080 5.420 1.240 ;
        RECT  5.020 0.470 5.140 1.240 ;
        RECT  3.280 0.470 5.020 0.590 ;
        RECT  3.120 0.470 3.280 1.710 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.050 ;
        LAYER M1 ;
        RECT  3.830 0.760 3.895 0.920 ;
        RECT  3.850 1.650 3.895 2.030 ;
        RECT  4.745 0.760 4.820 0.920 ;
        RECT  4.745 1.650 4.800 2.030 ;
        RECT  5.310 0.490 5.495 0.870 ;
        RECT  5.310 1.650 5.495 2.030 ;
    END
END LHCND4

MACRO LHCSND1
    CLASS CORE ;
    FOREIGN LHCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.080 2.970 1.240 ;
        RECT  2.970 1.005 3.110 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.600 3.930 1.760 ;
        RECT  3.790 0.760 3.930 0.920 ;
        RECT  3.930 0.760 4.070 1.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.940 4.540 2.100 ;
        RECT  4.540 1.390 4.590 2.100 ;
        RECT  4.540 0.420 4.590 0.955 ;
        RECT  4.590 0.420 4.710 2.100 ;
        RECT  4.710 1.940 4.730 2.100 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.395 1.320 1.520 ;
        RECT  1.320 0.860 1.480 1.520 ;
        RECT  1.480 1.360 2.110 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.015 1.050 1.235 ;
        RECT  1.050 0.725 1.190 1.235 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.015 0.730 1.235 ;
        RECT  0.730 0.725 0.870 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.550 3.390 2.050 ;
        RECT  1.650 1.650 2.330 1.810 ;
        RECT  1.400 0.570 2.330 0.730 ;
        RECT  2.330 0.570 2.450 1.810 ;
        RECT  2.450 1.080 2.670 1.240 ;
        RECT  0.220 1.440 0.260 2.050 ;
        RECT  0.220 0.610 0.260 0.850 ;
        RECT  0.260 1.930 1.490 2.050 ;
        RECT  1.490 1.930 1.730 2.090 ;
        RECT  2.900 0.550 3.230 0.710 ;
        RECT  2.870 1.930 3.230 2.050 ;
        RECT  2.710 1.700 2.870 2.050 ;
        RECT  2.340 1.930 2.710 2.050 ;
        RECT  4.390 1.050 4.460 1.270 ;
        RECT  4.270 1.050 4.390 2.000 ;
        RECT  3.660 1.880 4.270 2.000 ;
        RECT  3.660 0.420 3.800 0.580 ;
        RECT  3.520 0.420 3.660 2.000 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 1.650 1.810 ;
        RECT  0.100 0.610 0.220 2.050 ;
    END
END LHCSND1

MACRO LHCSND2
    CLASS CORE ;
    FOREIGN LHCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.960 3.130 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.960 4.090 2.100 ;
        RECT  4.090 1.390 4.250 2.100 ;
        RECT  4.040 0.710 4.250 0.870 ;
        RECT  4.250 1.960 4.280 2.100 ;
        RECT  4.250 0.710 4.390 1.525 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.780 1.940 4.810 2.100 ;
        RECT  4.810 1.390 4.890 2.100 ;
        RECT  4.810 0.420 4.890 0.900 ;
        RECT  4.890 0.420 4.970 2.100 ;
        RECT  4.970 1.940 5.000 2.100 ;
        RECT  4.970 0.780 5.030 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.395 1.320 1.520 ;
        RECT  1.320 0.860 1.480 1.520 ;
        RECT  1.480 1.360 2.110 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.015 1.050 1.235 ;
        RECT  1.050 0.725 1.190 1.235 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.015 0.730 1.235 ;
        RECT  0.730 0.725 0.870 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 2.330 0.300 ;
        RECT  2.330 -0.300 2.550 0.340 ;
        RECT  2.550 -0.300 3.660 0.300 ;
        RECT  3.660 -0.300 3.880 0.340 ;
        RECT  3.880 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 3.660 2.820 ;
        RECT  3.660 2.180 3.880 2.820 ;
        RECT  3.880 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.260 1.930 1.490 2.050 ;
        RECT  1.490 1.930 1.730 2.090 ;
        RECT  0.220 0.610 0.260 0.850 ;
        RECT  0.220 1.440 0.260 2.050 ;
        RECT  2.450 1.050 2.610 1.270 ;
        RECT  2.330 0.570 2.450 1.810 ;
        RECT  1.400 0.570 2.330 0.730 ;
        RECT  1.650 1.650 2.330 1.810 ;
        RECT  3.740 1.030 3.900 1.910 ;
        RECT  2.850 1.750 3.740 1.910 ;
        RECT  2.850 0.550 3.230 0.710 ;
        RECT  2.730 0.550 2.850 1.910 ;
        RECT  2.610 1.750 2.730 2.050 ;
        RECT  2.340 1.930 2.610 2.050 ;
        RECT  4.670 1.080 4.770 1.240 ;
        RECT  4.550 0.470 4.670 1.240 ;
        RECT  3.530 0.470 4.550 0.590 ;
        RECT  3.370 0.470 3.530 1.630 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 1.650 1.810 ;
        RECT  0.100 0.610 0.220 2.050 ;
    END
END LHCSND2

MACRO LHCSND4
    CLASS CORE ;
    FOREIGN LHCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.130 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.650 4.430 2.030 ;
        RECT  3.990 0.760 4.430 0.920 ;
        RECT  4.430 0.760 4.850 2.030 ;
        RECT  4.850 1.650 4.920 2.030 ;
        RECT  4.850 0.760 4.940 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 1.650 5.710 2.030 ;
        RECT  5.390 0.490 5.710 0.870 ;
        RECT  5.710 0.490 6.130 2.030 ;
        RECT  6.130 1.650 6.300 2.030 ;
        RECT  6.130 0.490 6.300 0.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.395 1.320 1.520 ;
        RECT  1.320 0.860 1.480 1.520 ;
        RECT  1.480 1.360 2.110 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.015 1.050 1.235 ;
        RECT  1.050 0.725 1.190 1.235 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.015 0.730 1.235 ;
        RECT  0.730 0.725 0.870 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 2.320 0.300 ;
        RECT  2.320 -0.300 2.540 0.340 ;
        RECT  2.540 -0.300 3.610 0.300 ;
        RECT  3.610 -0.300 3.830 0.340 ;
        RECT  3.830 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 3.610 2.820 ;
        RECT  3.610 2.180 3.830 2.820 ;
        RECT  3.830 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.490 1.930 1.730 2.090 ;
        RECT  0.260 1.930 1.490 2.050 ;
        RECT  0.220 0.610 0.260 0.850 ;
        RECT  0.220 1.440 0.260 2.050 ;
        RECT  2.450 1.050 2.610 1.270 ;
        RECT  2.330 0.570 2.450 1.810 ;
        RECT  1.400 0.570 2.330 0.730 ;
        RECT  1.650 1.650 2.330 1.810 ;
        RECT  3.730 1.030 3.890 1.910 ;
        RECT  2.850 1.750 3.730 1.910 ;
        RECT  2.850 0.550 3.210 0.710 ;
        RECT  2.730 0.550 2.850 1.910 ;
        RECT  2.610 1.750 2.730 2.050 ;
        RECT  2.340 1.930 2.610 2.050 ;
        RECT  5.270 1.080 5.495 1.240 ;
        RECT  5.150 0.470 5.270 1.240 ;
        RECT  3.510 0.470 5.150 0.590 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 1.650 1.810 ;
        RECT  3.350 0.470 3.510 1.630 ;
        RECT  0.100 0.610 0.220 2.050 ;
        LAYER M1 ;
        RECT  3.990 0.760 4.215 0.920 ;
        RECT  4.010 1.650 4.215 2.030 ;
        RECT  5.390 0.490 5.495 0.870 ;
        RECT  5.390 1.650 5.495 2.030 ;
    END
END LHCSND4

MACRO LHD1
    CLASS CORE ;
    FOREIGN LHD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.940 3.910 2.100 ;
        RECT  3.910 0.420 4.070 2.100 ;
        RECT  4.070 1.940 4.100 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.940 3.150 2.100 ;
        RECT  3.150 1.390 3.290 2.100 ;
        RECT  3.120 0.710 3.290 0.870 ;
        RECT  3.290 0.710 3.310 2.100 ;
        RECT  3.310 1.940 3.340 2.100 ;
        RECT  3.310 0.710 3.430 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.430 2.820 ;
        RECT  0.430 2.180 0.650 2.820 ;
        RECT  0.650 2.220 1.170 2.820 ;
        RECT  1.170 1.640 1.390 2.820 ;
        RECT  1.390 2.220 2.370 2.820 ;
        RECT  2.370 2.180 2.590 2.820 ;
        RECT  2.590 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.630 0.760 1.750 2.050 ;
        RECT  1.750 0.870 1.890 1.030 ;
        RECT  1.750 1.930 1.980 2.050 ;
        RECT  1.980 1.930 2.220 2.090 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  0.420 0.690 0.540 1.800 ;
        RECT  0.540 1.080 0.810 1.240 ;
        RECT  1.050 0.760 1.630 0.880 ;
        RECT  0.930 0.720 1.050 1.710 ;
        RECT  0.810 0.720 0.930 0.880 ;
        RECT  2.130 1.190 2.760 1.350 ;
        RECT  2.060 0.480 2.130 1.350 ;
        RECT  2.010 0.480 2.060 1.810 ;
        RECT  1.780 0.480 2.010 0.640 ;
        RECT  1.940 1.190 2.010 1.810 ;
        RECT  3.750 1.050 3.790 1.290 ;
        RECT  3.630 0.470 3.750 1.290 ;
        RECT  3.000 0.470 3.630 0.590 ;
        RECT  2.880 0.470 3.000 1.880 ;
        RECT  2.490 0.470 2.880 0.630 ;
        RECT  2.750 1.720 2.880 1.880 ;
        RECT  2.330 0.470 2.490 1.040 ;
        RECT  1.870 1.590 1.940 1.810 ;
        RECT  0.810 1.550 0.930 1.710 ;
        RECT  0.070 1.640 0.420 1.800 ;
    END
END LHD1

MACRO LHD2
    CLASS CORE ;
    FOREIGN LHD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.940 4.190 2.100 ;
        RECT  4.190 1.390 4.250 2.100 ;
        RECT  4.190 0.420 4.250 0.900 ;
        RECT  4.250 0.420 4.350 2.100 ;
        RECT  4.350 1.940 4.380 2.100 ;
        RECT  4.350 0.780 4.390 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.940 3.500 2.100 ;
        RECT  3.500 1.390 3.610 2.100 ;
        RECT  3.450 0.710 3.610 0.870 ;
        RECT  3.610 0.710 3.660 2.100 ;
        RECT  3.660 1.940 3.690 2.100 ;
        RECT  3.660 0.710 3.750 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.430 2.820 ;
        RECT  0.430 2.180 0.650 2.820 ;
        RECT  0.650 2.220 1.170 2.820 ;
        RECT  1.170 1.640 1.390 2.820 ;
        RECT  1.390 2.220 2.400 2.820 ;
        RECT  2.400 2.180 2.620 2.820 ;
        RECT  2.620 2.220 3.070 2.820 ;
        RECT  3.070 2.180 3.290 2.820 ;
        RECT  3.290 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.810 1.240 ;
        RECT  0.420 0.690 0.540 1.800 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  1.980 1.930 2.220 2.090 ;
        RECT  1.750 1.930 1.980 2.050 ;
        RECT  1.750 0.870 1.890 1.030 ;
        RECT  1.630 0.760 1.750 2.050 ;
        RECT  1.050 0.760 1.630 0.880 ;
        RECT  0.930 0.720 1.050 1.710 ;
        RECT  0.810 0.720 0.930 0.880 ;
        RECT  2.130 1.190 2.790 1.350 ;
        RECT  2.060 0.480 2.130 1.350 ;
        RECT  2.010 0.480 2.060 1.810 ;
        RECT  1.780 0.480 2.010 0.640 ;
        RECT  1.940 1.190 2.010 1.810 ;
        RECT  4.030 1.050 4.130 1.270 ;
        RECT  3.890 0.470 4.030 1.270 ;
        RECT  3.030 0.470 3.890 0.590 ;
        RECT  2.910 0.470 3.030 1.880 ;
        RECT  2.470 0.470 2.910 0.630 ;
        RECT  2.780 1.720 2.910 1.880 ;
        RECT  2.310 0.470 2.470 1.040 ;
        RECT  1.870 1.590 1.940 1.810 ;
        RECT  0.810 1.550 0.930 1.710 ;
        RECT  0.070 1.640 0.420 1.800 ;
    END
END LHD2

MACRO LHD4
    CLASS CORE ;
    FOREIGN LHD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.750 1.650 5.070 2.030 ;
        RECT  4.750 0.490 5.070 0.870 ;
        RECT  5.070 0.490 5.490 2.030 ;
        RECT  5.490 1.650 5.660 2.030 ;
        RECT  5.490 0.490 5.660 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.650 3.470 2.030 ;
        RECT  3.350 0.760 3.470 0.920 ;
        RECT  3.470 0.760 3.890 2.030 ;
        RECT  3.890 1.650 4.280 2.030 ;
        RECT  3.890 0.760 4.300 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.030 1.370 1.250 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.390 0.300 ;
        RECT  0.390 -0.300 0.610 0.340 ;
        RECT  0.610 -0.300 1.110 0.300 ;
        RECT  1.110 -0.300 1.330 0.340 ;
        RECT  1.330 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.390 2.820 ;
        RECT  0.390 2.180 0.610 2.820 ;
        RECT  0.610 2.220 1.070 2.820 ;
        RECT  1.070 1.980 1.290 2.820 ;
        RECT  1.290 2.220 2.320 2.820 ;
        RECT  2.320 2.180 2.540 2.820 ;
        RECT  2.540 2.220 2.970 2.820 ;
        RECT  2.970 2.180 3.190 2.820 ;
        RECT  3.190 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.080 0.780 1.240 ;
        RECT  0.420 0.690 0.540 1.800 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  1.940 1.930 2.180 2.090 ;
        RECT  1.660 1.930 1.940 2.050 ;
        RECT  1.660 0.760 1.820 1.080 ;
        RECT  1.020 0.760 1.660 0.880 ;
        RECT  1.540 1.640 1.660 2.050 ;
        RECT  1.020 1.640 1.540 1.760 ;
        RECT  1.010 0.760 1.020 1.760 ;
        RECT  0.900 0.720 1.010 1.760 ;
        RECT  0.770 0.720 0.900 0.880 ;
        RECT  2.090 1.190 2.790 1.350 ;
        RECT  2.000 0.480 2.090 1.350 ;
        RECT  1.970 0.480 2.000 1.780 ;
        RECT  1.740 0.480 1.970 0.640 ;
        RECT  1.880 1.190 1.970 1.780 ;
        RECT  4.575 1.080 4.855 1.240 ;
        RECT  4.455 0.470 4.575 1.240 ;
        RECT  3.030 0.470 4.455 0.590 ;
        RECT  2.910 0.470 3.030 1.880 ;
        RECT  2.430 0.470 2.910 0.630 ;
        RECT  2.700 1.720 2.910 1.880 ;
        RECT  1.780 1.620 1.880 1.780 ;
        RECT  2.270 0.470 2.430 1.040 ;
        RECT  0.770 1.600 0.900 1.760 ;
        RECT  0.070 1.640 0.420 1.800 ;
        LAYER M1 ;
        RECT  4.105 0.760 4.300 0.920 ;
        RECT  4.105 1.650 4.280 2.030 ;
        RECT  4.750 0.490 4.855 0.870 ;
        RECT  4.750 1.650 4.855 2.030 ;
    END
END LHD4

MACRO LHSND1
    CLASS CORE ;
    FOREIGN LHSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.725 2.790 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.940 3.500 2.100 ;
        RECT  3.500 1.390 3.610 2.100 ;
        RECT  3.470 0.710 3.610 0.870 ;
        RECT  3.610 0.710 3.660 2.100 ;
        RECT  3.660 1.940 3.690 2.100 ;
        RECT  3.660 0.710 3.750 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.955 4.230 2.100 ;
        RECT  4.230 1.390 4.250 2.100 ;
        RECT  4.230 0.420 4.250 0.900 ;
        RECT  4.250 0.420 4.390 2.100 ;
        RECT  4.390 1.960 4.420 2.100 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.400 1.050 1.520 ;
        RECT  1.050 0.770 1.210 1.520 ;
        RECT  1.210 1.360 1.620 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.235 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 2.820 0.300 ;
        RECT  2.820 -0.300 3.040 0.340 ;
        RECT  3.040 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 2.720 2.820 ;
        RECT  2.720 2.180 2.940 2.820 ;
        RECT  2.940 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.240 0.420 0.260 0.640 ;
        RECT  0.260 1.930 1.070 2.050 ;
        RECT  1.070 1.930 1.310 2.090 ;
        RECT  0.240 1.490 0.260 2.050 ;
        RECT  2.060 0.480 2.220 1.810 ;
        RECT  1.150 0.480 2.060 0.640 ;
        RECT  2.950 1.030 3.110 1.480 ;
        RECT  2.510 1.360 2.950 1.480 ;
        RECT  2.500 0.440 2.710 0.600 ;
        RECT  2.500 1.360 2.510 2.050 ;
        RECT  2.350 0.440 2.500 2.050 ;
        RECT  1.890 1.930 2.350 2.050 ;
        RECT  4.090 1.040 4.130 1.280 ;
        RECT  3.970 0.470 4.090 1.280 ;
        RECT  3.350 0.470 3.970 0.590 ;
        RECT  3.230 0.470 3.350 1.760 ;
        RECT  3.100 0.710 3.230 0.870 ;
        RECT  3.100 1.600 3.230 1.760 ;
        RECT  1.650 1.930 1.890 2.090 ;
        RECT  1.180 1.650 2.060 1.810 ;
        RECT  0.100 0.420 0.240 2.050 ;
    END
END LHSND1

MACRO LHSND2
    CLASS CORE ;
    FOREIGN LHSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.940 3.640 2.100 ;
        RECT  3.610 0.710 3.640 1.515 ;
        RECT  3.640 0.710 3.750 2.100 ;
        RECT  3.750 1.390 3.800 2.100 ;
        RECT  3.800 1.940 3.830 2.100 ;
        RECT  3.750 0.710 3.850 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.390 1.940 4.420 2.100 ;
        RECT  4.420 1.390 4.570 2.100 ;
        RECT  4.420 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.580 2.100 ;
        RECT  4.580 1.940 4.610 2.100 ;
        RECT  4.580 0.780 4.710 1.515 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.080 0.410 1.300 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.400 1.040 1.520 ;
        RECT  1.040 0.750 1.200 1.520 ;
        RECT  1.200 1.360 1.540 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 0.800 0.730 1.020 ;
        RECT  0.730 0.725 0.870 1.235 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.700 0.340 ;
        RECT  0.700 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 3.220 0.300 ;
        RECT  3.220 -0.300 3.440 0.340 ;
        RECT  3.440 -0.300 4.000 0.300 ;
        RECT  4.000 -0.300 4.220 0.340 ;
        RECT  4.220 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.340 ;
        RECT  5.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.220 2.820 ;
        RECT  3.220 2.180 3.440 2.820 ;
        RECT  3.440 2.220 4.000 2.820 ;
        RECT  4.000 2.180 4.220 2.820 ;
        RECT  4.220 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 1.930 1.230 2.090 ;
        RECT  0.260 1.930 0.990 2.050 ;
        RECT  0.220 0.420 0.260 0.640 ;
        RECT  0.220 1.490 0.260 2.050 ;
        RECT  2.080 1.050 2.180 1.270 ;
        RECT  1.960 0.510 2.080 1.790 ;
        RECT  1.360 0.510 1.960 0.630 ;
        RECT  1.100 1.650 1.960 1.790 ;
        RECT  3.260 1.030 3.430 2.050 ;
        RECT  2.420 1.930 3.260 2.050 ;
        RECT  2.420 0.490 2.690 0.650 ;
        RECT  2.300 0.490 2.420 2.050 ;
        RECT  2.200 1.475 2.300 2.050 ;
        RECT  1.830 1.930 2.200 2.050 ;
        RECT  4.110 0.470 4.270 1.290 ;
        RECT  3.115 0.470 4.110 0.590 ;
        RECT  2.975 0.470 3.115 1.800 ;
        RECT  2.830 0.710 2.975 0.870 ;
        RECT  1.590 1.930 1.830 2.090 ;
        RECT  1.140 0.490 1.360 0.630 ;
        RECT  2.810 1.640 2.975 1.800 ;
        RECT  0.100 0.420 0.220 2.050 ;
    END
END LHSND2

MACRO LHSND4
    CLASS CORE ;
    FOREIGN LHSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.650 3.790 2.030 ;
        RECT  3.590 0.760 3.790 0.920 ;
        RECT  3.790 0.760 4.210 2.030 ;
        RECT  4.210 1.650 4.540 2.030 ;
        RECT  4.210 0.760 4.560 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.030 1.650 5.390 2.030 ;
        RECT  5.030 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.960 2.030 ;
        RECT  5.810 0.490 5.960 0.870 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.080 0.410 1.300 ;
        RECT  0.410 1.005 0.550 1.520 ;
        RECT  0.550 1.400 1.040 1.520 ;
        RECT  1.040 0.750 1.200 1.520 ;
        RECT  1.200 1.360 1.540 1.520 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 0.800 0.730 1.020 ;
        RECT  0.730 0.725 0.870 1.235 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.700 0.340 ;
        RECT  0.700 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 3.220 0.300 ;
        RECT  3.220 -0.300 3.440 0.340 ;
        RECT  3.440 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.220 2.820 ;
        RECT  3.220 2.180 3.440 2.820 ;
        RECT  3.440 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 1.930 1.230 2.090 ;
        RECT  0.260 1.930 0.990 2.050 ;
        RECT  0.220 0.420 0.260 0.640 ;
        RECT  0.220 1.490 0.260 2.050 ;
        RECT  2.080 1.050 2.180 1.270 ;
        RECT  1.960 0.510 2.080 1.790 ;
        RECT  1.360 0.510 1.960 0.630 ;
        RECT  1.100 1.650 1.960 1.790 ;
        RECT  3.260 1.030 3.430 2.050 ;
        RECT  2.420 1.930 3.260 2.050 ;
        RECT  2.420 0.490 2.690 0.650 ;
        RECT  2.300 0.490 2.420 2.050 ;
        RECT  2.200 1.475 2.300 2.050 ;
        RECT  1.830 1.930 2.200 2.050 ;
        RECT  4.870 1.080 5.140 1.240 ;
        RECT  4.750 0.470 4.870 1.240 ;
        RECT  3.115 0.470 4.750 0.590 ;
        RECT  2.975 0.470 3.115 1.800 ;
        RECT  2.830 0.710 2.975 0.870 ;
        RECT  1.590 1.930 1.830 2.090 ;
        RECT  2.810 1.640 2.975 1.800 ;
        RECT  1.140 0.490 1.360 0.630 ;
        RECT  0.100 0.420 0.220 2.050 ;
        LAYER M1 ;
        RECT  4.425 0.760 4.560 0.920 ;
        RECT  4.425 1.650 4.540 2.030 ;
        RECT  5.030 0.490 5.175 0.870 ;
        RECT  5.030 1.650 5.175 2.030 ;
    END
END LHSND4

MACRO LNCND1
    CLASS CORE ;
    FOREIGN LNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.940 3.830 2.100 ;
        RECT  3.830 1.390 3.930 2.100 ;
        RECT  3.780 0.710 3.930 0.870 ;
        RECT  3.930 0.710 3.990 2.100 ;
        RECT  3.990 1.940 4.020 2.100 ;
        RECT  3.990 0.710 4.070 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.940 4.550 2.100 ;
        RECT  4.550 1.390 4.570 2.100 ;
        RECT  4.550 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.710 2.100 ;
        RECT  4.710 1.940 4.740 2.100 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.580 2.050 ;
        RECT  1.580 1.930 1.820 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 3.130 0.300 ;
        RECT  3.130 -0.300 3.350 0.340 ;
        RECT  3.350 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.130 2.820 ;
        RECT  3.130 2.180 3.350 2.820 ;
        RECT  3.350 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.450 1.080 2.750 1.240 ;
        RECT  0.260 0.765 1.310 0.885 ;
        RECT  1.310 0.765 1.430 1.090 ;
        RECT  1.430 0.930 1.970 1.090 ;
        RECT  1.970 0.930 2.130 1.540 ;
        RECT  2.330 0.650 2.450 1.810 ;
        RECT  1.690 0.650 2.330 0.770 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  1.550 0.530 1.690 0.770 ;
        RECT  2.990 1.050 3.360 1.270 ;
        RECT  2.870 0.480 2.990 2.050 ;
        RECT  2.750 0.480 2.870 0.640 ;
        RECT  2.770 1.630 2.870 2.050 ;
        RECT  2.400 1.930 2.770 2.050 ;
        RECT  4.420 1.050 4.450 1.290 ;
        RECT  4.300 0.470 4.420 1.290 ;
        RECT  3.640 0.470 4.300 0.590 ;
        RECT  3.480 0.470 3.640 1.830 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.030 ;
    END
END LNCND1

MACRO LNCND2
    CLASS CORE ;
    FOREIGN LNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.790 1.940 3.820 2.100 ;
        RECT  3.820 1.390 3.930 2.100 ;
        RECT  3.770 0.710 3.930 0.870 ;
        RECT  3.930 0.710 3.980 2.100 ;
        RECT  3.980 1.940 4.010 2.100 ;
        RECT  3.980 0.710 4.070 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.940 4.510 2.100 ;
        RECT  4.510 1.390 4.570 2.100 ;
        RECT  4.510 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.670 2.100 ;
        RECT  4.670 1.940 4.700 2.100 ;
        RECT  4.670 0.780 4.710 1.515 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.580 2.050 ;
        RECT  1.580 1.930 1.820 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 3.390 0.300 ;
        RECT  3.390 -0.300 3.610 0.340 ;
        RECT  3.610 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.390 2.820 ;
        RECT  3.390 2.180 3.610 2.820 ;
        RECT  3.610 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 0.930 2.130 1.540 ;
        RECT  1.430 0.930 1.970 1.090 ;
        RECT  1.310 0.765 1.430 1.090 ;
        RECT  0.260 0.765 1.310 0.885 ;
        RECT  2.450 1.080 2.720 1.240 ;
        RECT  2.330 0.650 2.450 1.810 ;
        RECT  1.690 0.650 2.330 0.770 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  1.550 0.530 1.690 0.770 ;
        RECT  3.470 1.030 3.630 2.050 ;
        RECT  2.960 1.930 3.470 2.050 ;
        RECT  2.840 0.470 2.960 2.050 ;
        RECT  2.720 0.470 2.840 0.630 ;
        RECT  2.740 1.630 2.840 2.050 ;
        RECT  2.400 1.930 2.740 2.050 ;
        RECT  4.360 1.050 4.430 1.270 ;
        RECT  4.220 0.470 4.360 1.270 ;
        RECT  3.280 0.470 4.220 0.590 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.030 ;
        RECT  3.120 0.470 3.280 1.710 ;
    END
END LNCND2

MACRO LNCND4
    CLASS CORE ;
    FOREIGN LNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.650 4.110 2.030 ;
        RECT  3.830 0.760 4.110 0.920 ;
        RECT  4.110 0.760 4.530 2.030 ;
        RECT  4.530 1.650 4.800 2.030 ;
        RECT  4.530 0.760 4.820 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.310 1.650 5.710 2.030 ;
        RECT  5.310 0.490 5.710 0.870 ;
        RECT  5.710 0.490 6.130 2.030 ;
        RECT  6.130 1.650 6.260 2.030 ;
        RECT  6.130 0.490 6.260 0.870 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.580 2.050 ;
        RECT  1.580 1.930 1.820 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 3.450 0.300 ;
        RECT  3.450 -0.300 3.670 0.340 ;
        RECT  3.670 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.120 2.820 ;
        RECT  1.120 2.180 1.340 2.820 ;
        RECT  1.340 2.220 3.450 2.820 ;
        RECT  3.450 2.180 3.670 2.820 ;
        RECT  3.670 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.970 0.930 2.130 1.540 ;
        RECT  1.430 0.930 1.970 1.090 ;
        RECT  1.310 0.765 1.430 1.090 ;
        RECT  0.260 0.765 1.310 0.885 ;
        RECT  2.450 1.080 2.720 1.240 ;
        RECT  2.330 0.650 2.450 1.810 ;
        RECT  1.690 0.650 2.330 0.770 ;
        RECT  1.930 1.690 2.330 1.810 ;
        RECT  1.710 1.670 1.930 1.810 ;
        RECT  0.940 1.690 1.710 1.810 ;
        RECT  1.550 0.530 1.690 0.770 ;
        RECT  3.455 1.030 3.615 2.050 ;
        RECT  2.960 1.930 3.455 2.050 ;
        RECT  2.840 0.470 2.960 2.050 ;
        RECT  2.720 0.470 2.840 0.630 ;
        RECT  2.740 1.630 2.840 2.050 ;
        RECT  2.400 1.930 2.740 2.050 ;
        RECT  5.140 1.080 5.420 1.240 ;
        RECT  5.020 0.470 5.140 1.240 ;
        RECT  3.280 0.470 5.020 0.590 ;
        RECT  3.120 0.470 3.280 1.710 ;
        RECT  2.160 1.930 2.400 2.090 ;
        RECT  0.700 1.670 0.940 1.810 ;
        RECT  0.100 0.570 0.260 2.030 ;
        LAYER M1 ;
        RECT  3.830 0.760 3.895 0.920 ;
        RECT  3.850 1.650 3.895 2.030 ;
        RECT  4.745 0.760 4.820 0.920 ;
        RECT  4.745 1.650 4.800 2.030 ;
        RECT  5.310 0.490 5.495 0.870 ;
        RECT  5.310 1.650 5.495 2.030 ;
    END
END LNCND4

MACRO LNCSND1
    CLASS CORE ;
    FOREIGN LNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.080 2.970 1.240 ;
        RECT  2.970 1.005 3.110 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.600 3.930 1.760 ;
        RECT  3.790 0.760 3.930 0.920 ;
        RECT  3.930 0.760 4.070 1.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.940 4.540 2.100 ;
        RECT  4.540 1.390 4.590 2.100 ;
        RECT  4.540 0.420 4.590 0.955 ;
        RECT  4.590 0.420 4.710 2.100 ;
        RECT  4.710 1.940 4.730 2.100 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.490 2.050 ;
        RECT  1.490 1.930 1.730 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.220 1.470 0.260 1.710 ;
        RECT  0.220 0.550 0.260 0.880 ;
        RECT  0.260 0.760 1.320 0.880 ;
        RECT  1.320 0.760 1.480 1.520 ;
        RECT  1.480 1.360 2.110 1.520 ;
        RECT  2.450 1.080 2.670 1.240 ;
        RECT  2.330 0.480 2.450 1.810 ;
        RECT  1.410 0.480 2.330 0.640 ;
        RECT  3.230 0.490 3.390 2.050 ;
        RECT  2.900 0.490 3.230 0.650 ;
        RECT  2.680 1.890 3.230 2.050 ;
        RECT  2.340 1.930 2.680 2.050 ;
        RECT  4.390 1.050 4.460 1.270 ;
        RECT  4.270 1.050 4.390 2.000 ;
        RECT  3.660 1.880 4.270 2.000 ;
        RECT  3.660 0.420 3.800 0.570 ;
        RECT  3.520 0.420 3.660 2.000 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 2.330 1.810 ;
        RECT  0.100 0.550 0.220 1.710 ;
    END
END LNCSND1

MACRO LNCSND2
    CLASS CORE ;
    FOREIGN LNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 0.960 3.130 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.960 4.090 2.100 ;
        RECT  4.090 1.390 4.250 2.100 ;
        RECT  4.040 0.710 4.250 0.870 ;
        RECT  4.250 1.960 4.280 2.100 ;
        RECT  4.250 0.710 4.390 1.525 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.780 1.940 4.810 2.100 ;
        RECT  4.810 1.390 4.890 2.100 ;
        RECT  4.810 0.420 4.890 0.900 ;
        RECT  4.890 0.420 4.970 2.100 ;
        RECT  4.970 1.940 5.000 2.100 ;
        RECT  4.970 0.780 5.030 1.515 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.490 2.050 ;
        RECT  1.490 1.930 1.730 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 2.330 0.300 ;
        RECT  2.330 -0.300 2.550 0.340 ;
        RECT  2.550 -0.300 3.660 0.300 ;
        RECT  3.660 -0.300 3.880 0.340 ;
        RECT  3.880 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 3.660 2.820 ;
        RECT  3.660 2.180 3.880 2.820 ;
        RECT  3.880 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.360 2.110 1.520 ;
        RECT  1.320 0.760 1.480 1.520 ;
        RECT  0.260 0.760 1.320 0.880 ;
        RECT  0.220 0.550 0.260 0.880 ;
        RECT  0.220 1.470 0.260 1.710 ;
        RECT  2.450 1.050 2.610 1.270 ;
        RECT  2.330 0.480 2.450 1.810 ;
        RECT  1.410 0.480 2.330 0.640 ;
        RECT  3.740 1.030 3.900 1.910 ;
        RECT  2.850 1.750 3.740 1.910 ;
        RECT  2.850 0.490 3.230 0.650 ;
        RECT  2.730 0.490 2.850 1.910 ;
        RECT  2.610 1.750 2.730 2.050 ;
        RECT  2.340 1.930 2.610 2.050 ;
        RECT  4.670 1.080 4.770 1.240 ;
        RECT  4.550 0.470 4.670 1.240 ;
        RECT  3.530 0.470 4.550 0.590 ;
        RECT  3.370 0.470 3.530 1.630 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 2.330 1.810 ;
        RECT  0.100 0.550 0.220 1.710 ;
    END
END LNCSND2

MACRO LNCSND4
    CLASS CORE ;
    FOREIGN LNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.130 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.650 4.430 2.030 ;
        RECT  3.990 0.760 4.430 0.920 ;
        RECT  4.430 0.760 4.850 2.030 ;
        RECT  4.850 1.650 4.920 2.030 ;
        RECT  4.850 0.760 4.940 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.390 1.650 5.710 2.030 ;
        RECT  5.390 0.490 5.710 0.870 ;
        RECT  5.710 0.490 6.130 2.030 ;
        RECT  6.130 1.650 6.300 2.030 ;
        RECT  6.130 0.490 6.300 0.870 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.490 2.050 ;
        RECT  1.490 1.930 1.730 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END D
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 2.330 0.300 ;
        RECT  2.330 -0.300 2.550 0.340 ;
        RECT  2.550 -0.300 3.610 0.300 ;
        RECT  3.610 -0.300 3.830 0.340 ;
        RECT  3.830 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.360 2.820 ;
        RECT  0.360 2.180 0.580 2.820 ;
        RECT  0.580 2.220 1.110 2.820 ;
        RECT  1.110 2.180 1.330 2.820 ;
        RECT  1.330 2.220 3.080 2.820 ;
        RECT  3.080 2.180 3.300 2.820 ;
        RECT  3.300 2.220 3.610 2.820 ;
        RECT  3.610 2.180 3.830 2.820 ;
        RECT  3.830 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.480 1.360 2.110 1.520 ;
        RECT  1.320 0.760 1.480 1.520 ;
        RECT  0.260 0.760 1.320 0.880 ;
        RECT  0.220 0.550 0.260 0.880 ;
        RECT  0.220 1.470 0.260 1.710 ;
        RECT  2.450 1.050 2.610 1.270 ;
        RECT  2.330 0.480 2.450 1.810 ;
        RECT  1.410 0.480 2.330 0.640 ;
        RECT  3.730 1.030 3.890 1.910 ;
        RECT  2.850 1.750 3.730 1.910 ;
        RECT  2.850 0.490 3.210 0.650 ;
        RECT  2.730 0.490 2.850 1.910 ;
        RECT  2.610 1.750 2.730 2.050 ;
        RECT  2.340 1.930 2.610 2.050 ;
        RECT  5.270 1.080 5.495 1.240 ;
        RECT  5.150 0.470 5.270 1.240 ;
        RECT  3.510 0.470 5.150 0.590 ;
        RECT  3.350 0.470 3.510 1.630 ;
        RECT  2.100 1.930 2.340 2.090 ;
        RECT  0.690 1.670 2.330 1.810 ;
        RECT  0.100 0.550 0.220 1.710 ;
        LAYER M1 ;
        RECT  3.990 0.760 4.215 0.920 ;
        RECT  4.010 1.650 4.215 2.030 ;
        RECT  5.390 0.490 5.495 0.870 ;
        RECT  5.390 1.650 5.495 2.030 ;
    END
END LNCSND4

MACRO LND1
    CLASS CORE ;
    FOREIGN LND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.880 1.940 3.910 2.100 ;
        RECT  3.910 0.420 4.070 2.100 ;
        RECT  4.070 1.940 4.100 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.120 1.940 3.150 2.100 ;
        RECT  3.150 1.390 3.290 2.100 ;
        RECT  3.120 0.710 3.290 0.870 ;
        RECT  3.290 0.710 3.310 2.100 ;
        RECT  3.310 1.940 3.340 2.100 ;
        RECT  3.310 0.710 3.430 1.515 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.430 2.820 ;
        RECT  0.430 2.180 0.650 2.820 ;
        RECT  0.650 2.220 1.260 2.820 ;
        RECT  1.170 1.640 1.260 1.800 ;
        RECT  1.260 1.640 1.390 2.820 ;
        RECT  1.390 2.220 2.370 2.820 ;
        RECT  2.370 2.180 2.590 2.820 ;
        RECT  2.590 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 1.190 2.010 1.810 ;
        RECT  1.780 0.480 2.010 0.640 ;
        RECT  2.010 0.480 2.060 1.810 ;
        RECT  2.060 0.480 2.130 1.350 ;
        RECT  2.130 1.190 2.760 1.350 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  0.420 0.480 0.540 1.800 ;
        RECT  0.540 1.080 0.810 1.240 ;
        RECT  0.540 0.480 1.350 0.600 ;
        RECT  1.350 0.480 1.470 0.880 ;
        RECT  1.470 0.760 1.630 0.880 ;
        RECT  1.630 0.760 1.750 2.050 ;
        RECT  1.750 0.870 1.890 1.030 ;
        RECT  1.750 1.930 1.980 2.050 ;
        RECT  1.980 1.930 2.220 2.090 ;
        RECT  0.920 1.550 0.930 2.080 ;
        RECT  0.810 0.720 0.930 0.880 ;
        RECT  0.930 0.720 1.050 2.080 ;
        RECT  1.050 1.920 1.140 2.080 ;
        RECT  3.750 1.050 3.790 1.290 ;
        RECT  3.630 0.470 3.750 1.290 ;
        RECT  3.000 0.470 3.630 0.590 ;
        RECT  2.880 0.470 3.000 1.880 ;
        RECT  2.490 0.470 2.880 0.630 ;
        RECT  2.750 1.720 2.880 1.880 ;
        RECT  2.330 0.470 2.490 1.040 ;
        RECT  1.870 1.590 1.940 1.810 ;
        RECT  0.070 1.640 0.420 1.800 ;
        RECT  0.810 1.550 0.920 1.710 ;
    END
END LND1

MACRO LND2
    CLASS CORE ;
    FOREIGN LND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.940 4.190 2.100 ;
        RECT  4.190 1.390 4.250 2.100 ;
        RECT  4.190 0.420 4.250 0.900 ;
        RECT  4.250 0.420 4.350 2.100 ;
        RECT  4.350 1.940 4.380 2.100 ;
        RECT  4.350 0.780 4.390 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.940 3.500 2.100 ;
        RECT  3.500 1.390 3.610 2.100 ;
        RECT  3.450 0.710 3.610 0.870 ;
        RECT  3.610 0.710 3.660 2.100 ;
        RECT  3.660 1.940 3.690 2.100 ;
        RECT  3.660 0.710 3.750 1.515 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.430 2.820 ;
        RECT  0.430 2.180 0.650 2.820 ;
        RECT  0.650 2.220 1.260 2.820 ;
        RECT  1.170 1.640 1.260 1.800 ;
        RECT  1.260 1.640 1.390 2.820 ;
        RECT  1.390 2.220 2.400 2.820 ;
        RECT  2.400 2.180 2.620 2.820 ;
        RECT  2.620 2.220 3.070 2.820 ;
        RECT  3.070 2.180 3.290 2.820 ;
        RECT  3.290 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.050 1.920 1.140 2.080 ;
        RECT  0.930 0.720 1.050 2.080 ;
        RECT  0.810 0.720 0.930 0.880 ;
        RECT  0.920 1.550 0.930 2.080 ;
        RECT  1.980 1.930 2.220 2.090 ;
        RECT  1.750 1.930 1.980 2.050 ;
        RECT  1.750 0.870 1.890 1.030 ;
        RECT  1.630 0.760 1.750 2.050 ;
        RECT  1.520 0.760 1.630 0.880 ;
        RECT  1.400 0.480 1.520 0.880 ;
        RECT  0.540 0.480 1.400 0.600 ;
        RECT  0.540 1.080 0.810 1.240 ;
        RECT  0.420 0.480 0.540 1.800 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  2.130 1.190 2.790 1.350 ;
        RECT  2.060 0.480 2.130 1.350 ;
        RECT  2.010 0.480 2.060 1.810 ;
        RECT  1.780 0.480 2.010 0.640 ;
        RECT  1.940 1.190 2.010 1.810 ;
        RECT  4.030 1.050 4.130 1.270 ;
        RECT  3.890 0.470 4.030 1.270 ;
        RECT  3.030 0.470 3.890 0.590 ;
        RECT  2.910 0.470 3.030 1.880 ;
        RECT  2.470 0.470 2.910 0.630 ;
        RECT  2.780 1.720 2.910 1.880 ;
        RECT  1.870 1.590 1.940 1.810 ;
        RECT  0.070 1.640 0.420 1.800 ;
        RECT  0.810 1.550 0.920 1.710 ;
        RECT  2.310 0.470 2.470 1.040 ;
    END
END LND2

MACRO LND4
    CLASS CORE ;
    FOREIGN LND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.970 1.650 5.390 2.030 ;
        RECT  4.970 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.930 2.030 ;
        RECT  5.810 0.490 5.930 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.490 1.650 3.790 2.030 ;
        RECT  3.490 0.760 3.790 0.920 ;
        RECT  3.790 0.760 4.210 2.030 ;
        RECT  4.210 1.650 4.450 2.030 ;
        RECT  4.210 0.760 4.470 0.920 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.725 1.510 1.250 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 1.150 0.300 ;
        RECT  1.150 -0.300 1.370 0.340 ;
        RECT  1.370 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 1.270 2.820 ;
        RECT  1.170 1.390 1.270 1.810 ;
        RECT  1.270 1.390 1.390 2.820 ;
        RECT  1.390 2.220 2.410 2.820 ;
        RECT  2.410 2.180 2.630 2.820 ;
        RECT  2.630 2.220 3.090 2.820 ;
        RECT  3.090 2.180 3.310 2.820 ;
        RECT  3.310 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.030 1.930 1.140 2.090 ;
        RECT  0.910 0.710 1.030 2.090 ;
        RECT  0.790 0.710 0.910 0.870 ;
        RECT  2.000 1.930 2.240 2.090 ;
        RECT  1.750 1.930 2.000 2.050 ;
        RECT  1.750 0.840 1.820 1.060 ;
        RECT  1.630 0.470 1.750 2.050 ;
        RECT  0.540 0.470 1.630 0.590 ;
        RECT  0.540 1.080 0.790 1.240 ;
        RECT  0.420 0.470 0.540 1.800 ;
        RECT  0.070 0.690 0.420 0.850 ;
        RECT  2.970 1.030 3.130 1.510 ;
        RECT  2.060 1.390 2.970 1.510 ;
        RECT  1.940 0.480 2.060 1.810 ;
        RECT  1.870 0.480 1.940 0.700 ;
        RECT  4.760 1.080 5.080 1.240 ;
        RECT  4.640 0.470 4.760 1.240 ;
        RECT  3.370 0.470 4.640 0.630 ;
        RECT  3.250 0.470 3.370 1.880 ;
        RECT  2.490 0.470 3.250 0.630 ;
        RECT  2.790 1.720 3.250 1.880 ;
        RECT  1.870 1.590 1.940 1.810 ;
        RECT  2.330 0.470 2.490 1.270 ;
        RECT  0.070 1.640 0.420 1.800 ;
        RECT  0.790 1.550 0.910 1.710 ;
        LAYER M1 ;
        RECT  3.490 0.760 3.575 0.920 ;
        RECT  3.490 1.650 3.575 2.030 ;
        RECT  4.425 0.760 4.470 0.920 ;
        RECT  4.425 1.650 4.450 2.030 ;
        RECT  4.970 0.490 5.175 0.870 ;
        RECT  4.970 1.650 5.175 2.030 ;
    END
END LND4

MACRO LNSND1
    CLASS CORE ;
    FOREIGN LNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.725 2.790 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.940 3.500 2.100 ;
        RECT  3.500 1.390 3.610 2.100 ;
        RECT  3.470 0.710 3.610 0.870 ;
        RECT  3.610 0.710 3.660 2.100 ;
        RECT  3.660 1.940 3.690 2.100 ;
        RECT  3.660 0.710 3.750 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.200 1.955 4.230 2.100 ;
        RECT  4.230 1.390 4.250 2.100 ;
        RECT  4.230 0.420 4.250 0.900 ;
        RECT  4.250 0.420 4.390 2.100 ;
        RECT  4.390 1.960 4.420 2.100 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.070 2.050 ;
        RECT  1.070 1.930 1.310 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.710 0.340 ;
        RECT  0.710 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 2.820 0.300 ;
        RECT  2.820 -0.300 3.040 0.340 ;
        RECT  3.040 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 2.720 2.820 ;
        RECT  2.720 2.180 2.940 2.820 ;
        RECT  2.940 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.240 1.490 0.260 1.730 ;
        RECT  0.240 0.420 0.260 0.885 ;
        RECT  0.260 0.765 1.050 0.885 ;
        RECT  1.050 0.765 1.210 1.520 ;
        RECT  1.210 1.360 1.620 1.520 ;
        RECT  2.060 0.480 2.220 1.810 ;
        RECT  1.130 0.480 2.060 0.640 ;
        RECT  2.950 1.030 3.110 1.480 ;
        RECT  2.510 1.360 2.950 1.480 ;
        RECT  2.500 0.440 2.710 0.600 ;
        RECT  2.500 1.360 2.510 2.050 ;
        RECT  2.350 0.440 2.500 2.050 ;
        RECT  1.890 1.930 2.350 2.050 ;
        RECT  4.090 1.040 4.130 1.280 ;
        RECT  3.970 0.470 4.090 1.280 ;
        RECT  3.350 0.470 3.970 0.590 ;
        RECT  3.230 0.470 3.350 1.760 ;
        RECT  3.100 0.710 3.230 0.870 ;
        RECT  1.650 1.930 1.890 2.090 ;
        RECT  1.180 1.650 2.060 1.810 ;
        RECT  3.100 1.600 3.230 1.760 ;
        RECT  0.100 0.420 0.240 1.730 ;
    END
END LNSND1

MACRO LNSND2
    CLASS CORE ;
    FOREIGN LNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.940 3.640 2.100 ;
        RECT  3.610 0.710 3.640 1.515 ;
        RECT  3.640 0.710 3.750 2.100 ;
        RECT  3.750 1.390 3.800 2.100 ;
        RECT  3.800 1.940 3.830 2.100 ;
        RECT  3.750 0.710 3.850 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.390 1.940 4.420 2.100 ;
        RECT  4.420 1.390 4.570 2.100 ;
        RECT  4.420 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.580 2.100 ;
        RECT  4.580 1.940 4.610 2.100 ;
        RECT  4.580 0.780 4.710 1.515 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 0.990 2.050 ;
        RECT  0.990 1.930 1.230 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.700 0.340 ;
        RECT  0.700 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 3.220 0.300 ;
        RECT  3.220 -0.300 3.440 0.340 ;
        RECT  3.440 -0.300 4.000 0.300 ;
        RECT  4.000 -0.300 4.220 0.340 ;
        RECT  4.220 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.340 ;
        RECT  5.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.220 2.820 ;
        RECT  3.220 2.180 3.440 2.820 ;
        RECT  3.440 2.220 4.000 2.820 ;
        RECT  4.000 2.180 4.220 2.820 ;
        RECT  4.220 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 1.360 1.540 1.520 ;
        RECT  1.040 0.750 1.200 1.520 ;
        RECT  0.260 0.750 1.040 0.870 ;
        RECT  0.220 0.420 0.260 0.870 ;
        RECT  0.220 1.490 0.260 1.730 ;
        RECT  2.080 1.050 2.180 1.270 ;
        RECT  1.960 0.510 2.080 1.790 ;
        RECT  1.360 0.510 1.960 0.630 ;
        RECT  1.100 1.650 1.960 1.790 ;
        RECT  3.260 1.030 3.430 2.050 ;
        RECT  2.420 1.930 3.260 2.050 ;
        RECT  2.420 0.490 2.690 0.650 ;
        RECT  2.300 0.490 2.420 2.050 ;
        RECT  2.200 1.475 2.300 2.050 ;
        RECT  1.830 1.930 2.200 2.050 ;
        RECT  4.110 0.470 4.270 1.290 ;
        RECT  3.115 0.470 4.110 0.590 ;
        RECT  2.975 0.470 3.115 1.800 ;
        RECT  2.830 0.710 2.975 0.870 ;
        RECT  2.810 1.640 2.975 1.800 ;
        RECT  1.590 1.930 1.830 2.090 ;
        RECT  1.120 0.490 1.360 0.630 ;
        RECT  0.100 0.420 0.220 1.730 ;
    END
END LNSND2

MACRO LNSND4
    CLASS CORE ;
    FOREIGN LNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.650 3.790 2.030 ;
        RECT  3.590 0.760 3.790 0.920 ;
        RECT  3.790 0.760 4.210 2.030 ;
        RECT  4.210 1.650 4.540 2.030 ;
        RECT  4.210 0.760 4.560 0.920 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.030 1.650 5.390 2.030 ;
        RECT  5.030 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.960 2.030 ;
        RECT  5.810 0.490 5.960 0.870 ;
        END
    END Q
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 2.050 ;
        RECT  0.550 1.930 0.990 2.050 ;
        RECT  0.990 1.930 1.230 2.090 ;
        END
    END EN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.700 0.340 ;
        RECT  0.700 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 3.220 0.300 ;
        RECT  3.220 -0.300 3.440 0.340 ;
        RECT  3.440 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.410 2.820 ;
        RECT  0.410 2.180 0.630 2.820 ;
        RECT  0.630 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.220 2.820 ;
        RECT  3.220 2.180 3.440 2.820 ;
        RECT  3.440 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.200 1.360 1.540 1.520 ;
        RECT  1.040 0.750 1.200 1.520 ;
        RECT  0.260 0.750 1.040 0.870 ;
        RECT  0.220 0.420 0.260 0.870 ;
        RECT  0.220 1.490 0.260 1.730 ;
        RECT  2.080 1.050 2.180 1.270 ;
        RECT  1.960 0.510 2.080 1.790 ;
        RECT  1.360 0.510 1.960 0.630 ;
        RECT  1.100 1.650 1.960 1.790 ;
        RECT  3.260 1.030 3.430 2.050 ;
        RECT  2.420 1.930 3.260 2.050 ;
        RECT  2.420 0.490 2.690 0.650 ;
        RECT  2.300 0.490 2.420 2.050 ;
        RECT  2.200 1.475 2.300 2.050 ;
        RECT  1.830 1.930 2.200 2.050 ;
        RECT  4.870 1.080 5.140 1.240 ;
        RECT  4.750 0.470 4.870 1.240 ;
        RECT  3.115 0.470 4.750 0.590 ;
        RECT  2.975 0.470 3.115 1.800 ;
        RECT  2.830 0.710 2.975 0.870 ;
        RECT  1.590 1.930 1.830 2.090 ;
        RECT  1.120 0.490 1.360 0.630 ;
        RECT  2.810 1.640 2.975 1.800 ;
        RECT  0.100 0.420 0.220 1.730 ;
        LAYER M1 ;
        RECT  4.425 0.760 4.560 0.920 ;
        RECT  4.425 1.650 4.540 2.030 ;
        RECT  5.030 0.490 5.175 0.870 ;
        RECT  5.030 1.650 5.175 2.030 ;
    END
END LNSND4

MACRO MAOI222D0
    CLASS CORE ;
    FOREIGN MAOI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.820 0.410 1.980 ;
        RECT  0.070 0.710 0.410 0.870 ;
        RECT  0.410 0.710 0.550 1.980 ;
        RECT  1.510 0.710 1.670 1.125 ;
        RECT  0.550 1.635 2.010 1.770 ;
        RECT  1.670 1.005 2.010 1.125 ;
        RECT  2.010 1.005 2.150 1.770 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.830 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.710 0.300 ;
        RECT  0.710 -0.300 0.930 0.870 ;
        RECT  0.930 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.700 2.820 ;
        RECT  0.700 1.910 0.920 2.820 ;
        RECT  0.920 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.290 0.470 1.890 0.590 ;
        RECT  1.890 0.470 2.050 0.880 ;
        RECT  1.100 1.890 2.160 2.050 ;
        RECT  1.130 0.470 1.290 0.880 ;
    END
END MAOI222D0

MACRO MAOI222D1
    CLASS CORE ;
    FOREIGN MAOI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 0.765 0.260 1.755 ;
        RECT  0.260 0.765 0.270 2.055 ;
        RECT  0.270 0.465 0.290 2.055 ;
        RECT  0.290 1.635 0.480 2.055 ;
        RECT  0.290 0.465 0.490 0.885 ;
        RECT  0.480 1.635 2.330 1.795 ;
        RECT  1.700 0.710 2.330 0.830 ;
        RECT  2.330 0.710 2.470 1.795 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.285 1.150 1.515 ;
        RECT  1.150 1.190 1.370 1.515 ;
        RECT  1.370 1.285 1.510 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.950 0.930 1.390 ;
        RECT  0.930 0.950 1.630 1.070 ;
        RECT  1.630 0.950 1.750 1.390 ;
        RECT  1.750 1.005 1.785 1.390 ;
        RECT  1.785 1.005 2.150 1.235 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        RECT  0.960 -0.300 1.180 0.830 ;
        RECT  1.180 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.930 2.820 ;
        RECT  0.930 2.180 1.150 2.820 ;
        RECT  1.150 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.470 2.340 0.590 ;
        RECT  1.320 1.915 2.340 2.050 ;
        RECT  1.370 0.470 1.530 0.830 ;
    END
END MAOI222D1

MACRO MAOI222D2
    CLASS CORE ;
    FOREIGN MAOI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.960 3.230 2.100 ;
        RECT  3.230 1.390 3.280 2.100 ;
        RECT  3.230 0.420 3.280 0.900 ;
        RECT  3.280 0.420 3.390 2.100 ;
        RECT  3.390 1.960 3.420 2.100 ;
        RECT  3.390 0.780 3.440 1.515 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.285 1.100 1.515 ;
        RECT  1.100 1.210 1.320 1.515 ;
        RECT  1.320 1.285 1.510 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.970 0.930 1.390 ;
        RECT  0.930 0.970 1.670 1.090 ;
        RECT  1.670 0.970 1.830 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.930 0.300 ;
        RECT  0.930 -0.300 1.150 0.610 ;
        RECT  1.150 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.940 2.820 ;
        RECT  0.940 2.180 1.160 2.820 ;
        RECT  1.160 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.570 1.915 2.120 2.050 ;
        RECT  2.120 1.915 2.340 2.080 ;
        RECT  2.270 1.080 2.840 1.240 ;
        RECT  2.150 0.730 2.270 1.795 ;
        RECT  0.440 0.730 2.150 0.850 ;
        RECT  1.710 1.635 2.150 1.795 ;
        RECT  0.290 1.640 0.490 2.060 ;
        RECT  0.290 0.460 0.440 0.880 ;
        RECT  0.270 0.460 0.290 2.060 ;
        RECT  0.220 0.460 0.270 1.760 ;
        RECT  2.970 0.780 3.110 1.510 ;
        RECT  2.660 0.780 2.970 0.900 ;
        RECT  2.660 1.390 2.970 1.510 ;
        RECT  2.660 1.960 2.690 2.100 ;
        RECT  2.500 0.420 2.660 0.900 ;
        RECT  2.500 1.390 2.660 2.100 ;
        RECT  2.470 1.960 2.500 2.100 ;
        RECT  0.170 0.760 0.220 1.760 ;
        RECT  1.320 0.470 2.350 0.610 ;
        RECT  1.350 1.635 1.570 2.050 ;
    END
END MAOI222D2

MACRO MAOI222D4
    CLASS CORE ;
    FOREIGN MAOI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.640 3.470 2.020 ;
        RECT  3.150 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 4.060 2.020 ;
        RECT  3.890 0.500 4.060 0.880 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.285 1.100 1.515 ;
        RECT  1.100 1.210 1.320 1.515 ;
        RECT  1.320 1.285 1.510 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.970 0.930 1.390 ;
        RECT  0.930 0.970 1.670 1.090 ;
        RECT  1.670 0.970 1.830 1.515 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.930 0.300 ;
        RECT  0.930 -0.300 1.150 0.610 ;
        RECT  1.150 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.940 2.820 ;
        RECT  0.940 2.180 1.160 2.820 ;
        RECT  1.160 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.120 1.915 2.340 2.080 ;
        RECT  1.570 1.915 2.120 2.050 ;
        RECT  2.270 1.080 2.790 1.240 ;
        RECT  2.150 0.730 2.270 1.795 ;
        RECT  0.440 0.730 2.150 0.850 ;
        RECT  1.710 1.635 2.150 1.795 ;
        RECT  0.290 1.640 0.490 2.060 ;
        RECT  0.290 0.460 0.440 0.880 ;
        RECT  0.270 0.460 0.290 2.060 ;
        RECT  0.220 0.460 0.270 1.760 ;
        RECT  3.030 1.080 3.255 1.240 ;
        RECT  2.910 0.780 3.030 1.510 ;
        RECT  2.650 0.780 2.910 0.900 ;
        RECT  2.650 1.390 2.910 1.510 ;
        RECT  2.650 1.960 2.680 2.100 ;
        RECT  2.490 0.420 2.650 0.900 ;
        RECT  2.490 1.390 2.650 2.100 ;
        RECT  0.170 0.760 0.220 1.760 ;
        RECT  1.320 0.470 2.350 0.610 ;
        RECT  1.350 1.635 1.570 2.050 ;
        RECT  2.460 1.960 2.490 2.100 ;
        LAYER M1 ;
        RECT  3.150 1.640 3.255 2.020 ;
        RECT  3.150 0.500 3.255 0.880 ;
    END
END MAOI222D4

MACRO MAOI22D0
    CLASS CORE ;
    FOREIGN MAOI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 0.440 1.300 0.600 ;
        RECT  1.300 0.470 1.370 0.600 ;
        RECT  1.360 1.565 1.440 1.795 ;
        RECT  1.370 0.470 1.440 0.955 ;
        RECT  1.440 0.470 1.560 1.795 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.235 ;
        RECT  0.550 0.770 0.670 0.990 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 0.725 1.840 1.255 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.565 1.090 1.795 ;
        RECT  1.050 0.725 1.090 0.955 ;
        RECT  1.090 0.725 1.210 1.795 ;
        RECT  1.210 1.090 1.320 1.320 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.610 2.820 ;
        RECT  0.610 2.090 0.830 2.820 ;
        RECT  0.830 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.910 1.130 0.970 1.350 ;
        RECT  0.790 0.470 0.910 1.800 ;
        RECT  0.600 0.470 0.790 0.600 ;
        RECT  0.060 1.640 0.790 1.800 ;
        RECT  0.360 0.440 0.600 0.600 ;
    END
END MAOI22D0

MACRO MAOI22D1
    CLASS CORE ;
    FOREIGN MAOI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.180 0.430 1.400 0.850 ;
        RECT  1.530 1.635 2.010 1.795 ;
        RECT  1.400 0.725 2.010 0.850 ;
        RECT  2.010 0.725 2.150 1.795 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.080 0.790 1.240 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.840 0.300 ;
        RECT  1.840 -0.300 2.060 0.340 ;
        RECT  2.060 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.760 2.820 ;
        RECT  0.760 2.180 0.980 2.820 ;
        RECT  0.980 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.670 0.730 0.910 0.850 ;
        RECT  0.910 0.730 1.030 1.770 ;
        RECT  1.030 1.080 1.190 1.240 ;
        RECT  0.310 1.650 0.910 1.770 ;
        RECT  0.450 0.430 0.670 0.850 ;
        RECT  1.930 1.915 2.170 2.075 ;
        RECT  1.390 1.915 1.930 2.050 ;
        RECT  1.170 1.650 1.390 2.070 ;
        RECT  0.090 1.650 0.310 2.070 ;
    END
END MAOI22D1

MACRO MAOI22D2
    CLASS CORE ;
    FOREIGN MAOI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.960 2.550 2.100 ;
        RECT  2.550 1.390 2.650 2.100 ;
        RECT  2.550 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.710 2.100 ;
        RECT  2.710 1.960 2.740 2.100 ;
        RECT  2.710 0.780 2.790 1.515 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.700 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 1.080 1.150 1.240 ;
        RECT  0.820 0.765 0.940 1.770 ;
        RECT  0.280 0.765 0.820 0.885 ;
        RECT  0.660 1.650 0.820 1.770 ;
        RECT  0.440 1.650 0.660 2.070 ;
        RECT  1.830 0.450 2.070 0.610 ;
        RECT  1.290 0.490 1.830 0.610 ;
        RECT  2.270 0.730 2.430 1.755 ;
        RECT  1.430 0.730 2.270 0.885 ;
        RECT  1.400 1.635 2.270 1.755 ;
        RECT  1.180 1.635 1.400 2.050 ;
        RECT  1.070 0.470 1.290 0.890 ;
        RECT  0.060 0.470 0.280 0.885 ;
    END
END MAOI22D2

MACRO MAOI22D4
    CLASS CORE ;
    FOREIGN MAOI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.640 2.830 2.020 ;
        RECT  2.490 0.500 2.830 0.880 ;
        RECT  2.830 0.500 3.250 2.020 ;
        RECT  3.250 1.640 3.410 2.020 ;
        RECT  3.250 0.500 3.410 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.700 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 1.080 1.150 1.240 ;
        RECT  0.820 0.765 0.940 1.770 ;
        RECT  0.280 0.765 0.820 0.885 ;
        RECT  0.660 1.650 0.820 1.770 ;
        RECT  0.440 1.650 0.660 2.070 ;
        RECT  1.830 0.450 2.070 0.610 ;
        RECT  1.290 0.490 1.830 0.610 ;
        RECT  2.210 0.730 2.370 1.755 ;
        RECT  1.430 0.730 2.210 0.885 ;
        RECT  1.400 1.635 2.210 1.755 ;
        RECT  1.180 1.635 1.400 2.050 ;
        RECT  1.070 0.470 1.290 0.890 ;
        RECT  0.060 0.470 0.280 0.885 ;
        LAYER M1 ;
        RECT  2.490 0.500 2.615 0.880 ;
        RECT  2.490 1.640 2.615 2.020 ;
    END
END MAOI22D4

MACRO MOAI22D0
    CLASS CORE ;
    FOREIGN MOAI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.830 1.690 1.990 ;
        RECT  1.530 0.710 1.690 0.870 ;
        RECT  1.690 0.710 1.830 1.990 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.215 1.570 1.435 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.245 0.810 1.405 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.760 0.300 ;
        RECT  0.760 -0.300 0.980 0.340 ;
        RECT  0.980 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.870 2.820 ;
        RECT  0.870 2.180 1.090 2.820 ;
        RECT  1.090 2.220 1.900 2.820 ;
        RECT  1.900 2.180 2.120 2.820 ;
        RECT  2.120 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.080 1.245 1.240 1.405 ;
        RECT  0.960 0.710 1.080 1.990 ;
        RECT  0.070 0.710 0.960 0.870 ;
        RECT  1.960 0.470 2.120 0.880 ;
        RECT  1.360 0.470 1.960 0.590 ;
        RECT  1.200 0.470 1.360 0.880 ;
        RECT  0.460 1.830 0.960 1.990 ;
    END
END MOAI22D0

MACRO MOAI22D1
    CLASS CORE ;
    FOREIGN MOAI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.640 1.480 2.060 ;
        RECT  1.480 1.640 1.690 1.760 ;
        RECT  1.530 0.710 1.690 0.870 ;
        RECT  1.690 0.710 1.830 1.760 ;
        END
    END ZN
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.570 1.270 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.080 0.810 1.240 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.760 0.300 ;
        RECT  0.760 -0.300 0.980 0.340 ;
        RECT  0.980 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.870 2.820 ;
        RECT  0.870 2.180 1.090 2.820 ;
        RECT  1.090 2.220 1.900 2.820 ;
        RECT  1.900 2.180 2.120 2.820 ;
        RECT  2.120 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.310 0.690 0.930 0.850 ;
        RECT  0.930 0.690 1.050 1.760 ;
        RECT  1.050 1.075 1.250 1.235 ;
        RECT  0.700 1.640 0.930 1.760 ;
        RECT  0.480 1.640 0.700 2.060 ;
        RECT  2.120 0.430 2.150 0.570 ;
        RECT  1.960 0.430 2.120 0.880 ;
        RECT  1.930 0.430 1.960 0.590 ;
        RECT  1.390 0.470 1.930 0.590 ;
        RECT  0.090 0.430 0.310 0.850 ;
        RECT  1.170 0.470 1.390 0.880 ;
    END
END MOAI22D1

MACRO MOAI22D2
    CLASS CORE ;
    FOREIGN MOAI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.960 2.550 2.100 ;
        RECT  2.550 1.390 2.650 2.100 ;
        RECT  2.550 0.420 2.650 0.910 ;
        RECT  2.650 0.420 2.710 2.100 ;
        RECT  2.710 1.960 2.740 2.100 ;
        RECT  2.710 0.790 2.790 1.515 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.700 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 1.080 1.150 1.240 ;
        RECT  0.820 0.750 0.940 1.755 ;
        RECT  0.660 0.750 0.820 0.870 ;
        RECT  0.280 1.635 0.820 1.755 ;
        RECT  0.440 0.450 0.660 0.870 ;
        RECT  1.830 1.910 2.070 2.070 ;
        RECT  1.290 1.910 1.830 2.030 ;
        RECT  2.270 0.765 2.430 1.790 ;
        RECT  1.400 0.765 2.270 0.885 ;
        RECT  1.430 1.635 2.270 1.790 ;
        RECT  1.180 0.470 1.400 0.885 ;
        RECT  1.070 1.630 1.290 2.050 ;
        RECT  0.060 1.635 0.280 2.050 ;
    END
END MOAI22D2

MACRO MOAI22D4
    CLASS CORE ;
    FOREIGN MOAI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.640 2.830 2.020 ;
        RECT  2.490 0.500 2.830 0.880 ;
        RECT  2.830 0.500 3.250 2.020 ;
        RECT  3.250 1.640 3.410 2.020 ;
        RECT  3.250 0.500 3.410 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.700 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.940 1.080 1.150 1.240 ;
        RECT  0.820 0.750 0.940 1.755 ;
        RECT  0.660 0.750 0.820 0.870 ;
        RECT  0.280 1.635 0.820 1.755 ;
        RECT  0.440 0.450 0.660 0.870 ;
        RECT  1.830 1.910 2.070 2.070 ;
        RECT  1.290 1.910 1.830 2.030 ;
        RECT  2.210 0.765 2.370 1.790 ;
        RECT  1.400 0.765 2.210 0.885 ;
        RECT  1.430 1.635 2.210 1.790 ;
        RECT  1.180 0.470 1.400 0.885 ;
        RECT  1.070 1.630 1.290 2.050 ;
        RECT  0.060 1.635 0.280 2.050 ;
        LAYER M1 ;
        RECT  2.490 0.500 2.615 0.880 ;
        RECT  2.490 1.640 2.615 2.020 ;
    END
END MOAI22D4

MACRO MUX2D0
    CLASS CORE ;
    FOREIGN MUX2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.490 2.790 1.890 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.180 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.005 0.930 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.620 0.300 ;
        RECT  0.620 -0.300 0.780 0.800 ;
        RECT  0.780 -0.300 2.190 0.300 ;
        RECT  2.190 -0.300 2.410 0.340 ;
        RECT  2.410 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.580 2.820 ;
        RECT  0.580 1.920 0.800 2.820 ;
        RECT  0.800 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.470 2.510 1.290 ;
        RECT  1.870 0.710 1.990 0.870 ;
        RECT  1.870 1.640 2.010 1.800 ;
        RECT  0.190 0.590 0.370 0.750 ;
        RECT  0.370 0.590 0.490 1.800 ;
        RECT  0.490 1.680 0.965 1.800 ;
        RECT  0.965 1.680 1.085 2.040 ;
        RECT  1.085 1.920 1.520 2.040 ;
        RECT  1.520 1.920 1.760 2.080 ;
        RECT  0.950 0.590 1.090 0.750 ;
        RECT  1.090 0.590 1.210 1.560 ;
        RECT  1.580 0.470 2.350 0.590 ;
        RECT  1.420 0.470 1.580 1.790 ;
        RECT  1.750 0.710 1.870 1.800 ;
        RECT  1.330 0.590 1.420 0.750 ;
        RECT  0.170 1.640 0.370 1.800 ;
        RECT  0.990 1.400 1.090 1.560 ;
    END
END MUX2D0

MACRO MUX2D1
    CLASS CORE ;
    FOREIGN MUX2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.640 ;
        RECT  0.760 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.940 0.670 2.820 ;
        RECT  0.670 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.340 0.470 2.460 1.290 ;
        RECT  2.460 1.050 2.510 1.290 ;
        RECT  1.890 0.710 2.000 0.870 ;
        RECT  1.890 1.640 2.020 1.800 ;
        RECT  0.060 1.660 0.380 1.820 ;
        RECT  0.350 0.760 0.380 0.880 ;
        RECT  0.380 0.760 0.500 1.820 ;
        RECT  0.500 1.700 0.790 1.820 ;
        RECT  0.790 1.700 0.910 2.040 ;
        RECT  0.910 1.920 1.510 2.040 ;
        RECT  1.510 1.920 1.750 2.080 ;
        RECT  1.030 0.640 1.190 1.760 ;
        RECT  1.570 0.470 2.340 0.590 ;
        RECT  1.410 0.470 1.570 1.760 ;
        RECT  1.760 0.710 1.890 1.800 ;
        RECT  0.190 0.440 0.350 0.880 ;
        RECT  0.920 0.640 1.030 0.800 ;
        RECT  1.320 0.470 1.410 0.630 ;
    END
END MUX2D1

MACRO MUX2D2
    CLASS CORE ;
    FOREIGN MUX2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.960 2.550 2.100 ;
        RECT  2.550 1.390 2.650 2.100 ;
        RECT  2.550 0.420 2.650 0.910 ;
        RECT  2.650 0.420 2.710 2.100 ;
        RECT  2.710 1.960 2.740 2.100 ;
        RECT  2.710 0.790 2.790 1.515 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.640 ;
        RECT  0.760 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.940 0.670 2.820 ;
        RECT  0.670 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.510 1.920 1.750 2.080 ;
        RECT  1.030 0.640 1.190 1.760 ;
        RECT  0.910 1.920 1.510 2.040 ;
        RECT  0.790 1.700 0.910 2.040 ;
        RECT  0.500 1.700 0.790 1.820 ;
        RECT  0.380 0.760 0.500 1.820 ;
        RECT  0.350 0.760 0.380 0.880 ;
        RECT  0.060 1.660 0.380 1.820 ;
        RECT  1.890 1.640 2.020 1.800 ;
        RECT  1.890 0.710 2.000 0.870 ;
        RECT  2.430 1.080 2.530 1.240 ;
        RECT  2.310 0.470 2.430 1.240 ;
        RECT  1.570 0.470 2.310 0.590 ;
        RECT  1.410 0.470 1.570 1.760 ;
        RECT  1.760 0.710 1.890 1.800 ;
        RECT  0.190 0.440 0.350 0.880 ;
        RECT  0.920 0.640 1.030 0.800 ;
        RECT  1.320 0.470 1.410 0.630 ;
    END
END MUX2D2

MACRO MUX2D4
    CLASS CORE ;
    FOREIGN MUX2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.650 3.790 2.030 ;
        RECT  3.470 0.490 3.790 0.870 ;
        RECT  3.790 0.490 4.210 2.030 ;
        RECT  4.210 1.650 4.380 2.030 ;
        RECT  4.210 0.490 4.380 0.870 ;
        END
    END Z
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.005 2.480 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.005 3.110 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.560 0.300 ;
        RECT  0.560 -0.300 0.780 0.340 ;
        RECT  0.780 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.970 0.430 1.190 0.850 ;
        RECT  0.900 1.390 1.060 1.930 ;
        RECT  0.360 0.690 0.970 0.850 ;
        RECT  0.260 1.390 0.900 1.510 ;
        RECT  0.260 0.430 0.360 0.850 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.140 0.430 0.260 2.100 ;
        RECT  0.100 1.390 0.140 2.100 ;
        RECT  2.200 1.650 2.330 1.810 ;
        RECT  2.200 0.710 2.320 0.870 ;
        RECT  2.080 0.710 2.200 1.810 ;
        RECT  2.810 0.710 3.020 0.870 ;
        RECT  2.810 1.890 3.020 2.050 ;
        RECT  2.690 0.710 2.810 2.050 ;
        RECT  1.860 1.930 2.690 2.050 ;
        RECT  1.810 0.710 1.960 0.870 ;
        RECT  1.810 1.410 1.860 2.050 ;
        RECT  1.700 0.710 1.810 2.050 ;
        RECT  3.350 1.080 3.575 1.240 ;
        RECT  3.230 0.470 3.350 1.240 ;
        RECT  1.570 0.470 3.230 0.590 ;
        RECT  1.480 0.470 1.570 0.630 ;
        RECT  1.690 0.710 1.700 1.530 ;
        RECT  1.320 0.470 1.480 1.910 ;
        RECT  1.930 1.100 2.080 1.260 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  3.470 1.650 3.575 2.030 ;
        RECT  3.470 0.490 3.575 0.870 ;
    END
END MUX2D4

MACRO MUX2ND0
    CLASS CORE ;
    FOREIGN MUX2ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 0.710 1.200 1.660 ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.770 0.420 1.010 0.590 ;
        RECT  1.010 0.470 2.010 0.590 ;
        RECT  2.010 0.470 2.070 1.515 ;
        RECT  2.070 0.420 2.150 1.515 ;
        RECT  2.150 0.420 2.330 0.560 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.810 2.820 ;
        RECT  1.810 1.970 2.030 2.820 ;
        RECT  2.030 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.710 2.430 1.850 ;
        RECT  1.690 1.730 2.270 1.850 ;
        RECT  1.570 1.730 1.690 2.050 ;
        RECT  1.010 1.930 1.570 2.050 ;
        RECT  1.430 0.710 1.570 1.610 ;
        RECT  0.770 1.930 1.010 2.090 ;
        RECT  0.570 0.710 0.730 1.660 ;
    END
END MUX2ND0

MACRO MUX2ND1
    CLASS CORE ;
    FOREIGN MUX2ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.960 3.270 2.100 ;
        RECT  3.270 0.420 3.430 2.100 ;
        RECT  3.430 1.960 3.460 2.100 ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.270 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.600 ;
        RECT  0.760 -0.300 2.140 0.300 ;
        RECT  2.140 -0.300 2.360 0.340 ;
        RECT  2.360 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.040 2.820 ;
        RECT  2.040 2.180 2.260 2.820 ;
        RECT  2.260 2.220 2.830 2.820 ;
        RECT  2.830 2.180 3.050 2.820 ;
        RECT  3.050 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.930 1.910 1.360 2.050 ;
        RECT  1.360 1.910 1.600 2.070 ;
        RECT  0.990 0.630 1.130 1.560 ;
        RECT  0.810 1.680 0.930 2.050 ;
        RECT  0.260 1.680 0.810 1.800 ;
        RECT  0.260 0.710 0.380 0.870 ;
        RECT  1.820 0.730 1.970 0.890 ;
        RECT  2.690 0.820 2.850 1.270 ;
        RECT  2.390 0.820 2.690 0.940 ;
        RECT  2.270 0.470 2.390 0.940 ;
        RECT  1.560 0.470 2.270 0.610 ;
        RECT  1.440 0.470 1.560 0.630 ;
        RECT  3.020 0.470 3.150 1.660 ;
        RECT  2.510 0.470 3.020 0.630 ;
        RECT  1.280 0.470 1.440 1.760 ;
        RECT  1.660 0.730 1.820 1.760 ;
        RECT  0.100 0.710 0.260 1.800 ;
        RECT  0.850 1.400 0.990 1.560 ;
        RECT  2.400 1.500 3.020 1.660 ;
    END
END MUX2ND1

MACRO MUX2ND2
    CLASS CORE ;
    FOREIGN MUX2ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.200 1.960 3.230 2.100 ;
        RECT  3.230 1.390 3.290 2.100 ;
        RECT  3.230 0.420 3.290 0.900 ;
        RECT  3.290 0.420 3.390 2.100 ;
        RECT  3.390 1.960 3.420 2.100 ;
        RECT  3.390 0.780 3.430 1.515 ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.725 0.870 1.270 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.540 0.300 ;
        RECT  0.540 -0.300 0.760 0.600 ;
        RECT  0.760 -0.300 2.140 0.300 ;
        RECT  2.140 -0.300 2.360 0.340 ;
        RECT  2.360 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.040 2.820 ;
        RECT  2.040 2.180 2.260 2.820 ;
        RECT  2.260 2.220 2.810 2.820 ;
        RECT  2.810 2.180 3.030 2.820 ;
        RECT  3.030 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.630 1.130 1.560 ;
        RECT  1.360 1.910 1.600 2.070 ;
        RECT  0.930 1.910 1.360 2.050 ;
        RECT  0.810 1.680 0.930 2.050 ;
        RECT  0.260 1.680 0.810 1.800 ;
        RECT  0.260 0.710 0.380 0.870 ;
        RECT  1.820 0.730 1.970 0.890 ;
        RECT  2.690 0.820 2.850 1.270 ;
        RECT  2.390 0.820 2.690 0.940 ;
        RECT  2.270 0.470 2.390 0.940 ;
        RECT  1.560 0.470 2.270 0.610 ;
        RECT  1.440 0.470 1.560 0.630 ;
        RECT  3.110 1.050 3.170 1.270 ;
        RECT  2.990 0.470 3.110 1.660 ;
        RECT  2.510 0.470 2.990 0.630 ;
        RECT  1.280 0.470 1.440 1.760 ;
        RECT  1.660 0.730 1.820 1.760 ;
        RECT  2.400 1.500 2.990 1.660 ;
        RECT  0.100 0.710 0.260 1.800 ;
        RECT  0.850 1.400 0.990 1.560 ;
    END
END MUX2ND2

MACRO MUX2ND4
    CLASS CORE ;
    FOREIGN MUX2ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.650 4.750 2.030 ;
        RECT  4.430 0.490 4.750 0.870 ;
        RECT  4.750 0.490 5.170 2.030 ;
        RECT  5.170 1.650 5.340 2.030 ;
        RECT  5.170 0.490 5.340 0.870 ;
        END
    END ZN
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.570 ;
        RECT  0.680 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.570 ;
        RECT  1.470 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 1.240 2.820 ;
        RECT  1.240 2.030 1.460 2.820 ;
        RECT  1.460 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.730 0.690 1.850 1.610 ;
        RECT  0.830 0.690 1.730 0.850 ;
        RECT  2.150 1.930 2.390 2.100 ;
        RECT  1.805 1.930 2.150 2.050 ;
        RECT  1.685 1.730 1.805 2.050 ;
        RECT  0.510 1.730 1.685 1.870 ;
        RECT  0.390 0.700 0.510 1.870 ;
        RECT  0.070 0.700 0.390 0.860 ;
        RECT  3.230 0.470 3.350 1.550 ;
        RECT  3.100 0.470 3.230 0.885 ;
        RECT  2.360 1.410 3.230 1.550 ;
        RECT  3.730 1.030 3.890 1.790 ;
        RECT  2.160 1.670 3.730 1.790 ;
        RECT  2.160 0.640 2.250 0.800 ;
        RECT  4.310 1.080 4.535 1.240 ;
        RECT  4.170 0.710 4.310 2.050 ;
        RECT  3.960 0.710 4.170 0.870 ;
        RECT  3.720 1.910 4.170 2.050 ;
        RECT  2.000 0.640 2.160 1.790 ;
        RECT  2.390 0.470 3.100 0.630 ;
        RECT  0.070 1.710 0.390 1.870 ;
        RECT  0.830 1.450 1.730 1.610 ;
        RECT  3.740 0.450 3.960 0.870 ;
        LAYER M1 ;
        RECT  4.430 0.490 4.535 0.870 ;
        RECT  4.430 1.650 4.535 2.030 ;
    END
END MUX2ND4

MACRO MUX3D0
    CLASS CORE ;
    FOREIGN MUX3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.470 1.770 4.570 1.930 ;
        RECT  4.470 0.710 4.570 0.870 ;
        RECT  4.570 0.710 4.710 1.930 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.490 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 0.985 0.410 1.225 ;
        RECT  0.410 0.985 0.550 1.515 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 0.890 1.250 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.590 0.300 ;
        RECT  0.590 -0.300 0.810 0.600 ;
        RECT  0.810 -0.300 2.170 0.300 ;
        RECT  2.170 -0.300 2.390 0.340 ;
        RECT  2.390 -0.300 4.100 0.300 ;
        RECT  4.100 -0.300 4.320 0.340 ;
        RECT  4.320 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.500 2.820 ;
        RECT  0.500 2.000 0.720 2.820 ;
        RECT  0.720 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.560 0.470 2.960 0.590 ;
        RECT  2.960 0.470 3.120 1.910 ;
        RECT  2.550 0.710 2.700 0.870 ;
        RECT  2.700 0.710 2.840 1.670 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.710 2.010 0.870 ;
        RECT  0.250 1.450 0.290 1.880 ;
        RECT  0.250 0.590 0.430 0.750 ;
        RECT  0.290 1.760 0.965 1.880 ;
        RECT  0.965 1.760 1.085 2.050 ;
        RECT  1.085 1.910 1.500 2.050 ;
        RECT  1.500 1.910 1.720 2.070 ;
        RECT  1.020 0.540 1.180 1.640 ;
        RECT  3.810 0.720 3.940 0.880 ;
        RECT  3.810 1.700 3.930 1.860 ;
        RECT  4.350 1.210 4.450 1.370 ;
        RECT  4.230 0.480 4.350 1.370 ;
        RECT  3.500 0.480 4.230 0.600 ;
        RECT  3.690 0.720 3.810 1.860 ;
        RECT  1.400 0.470 1.560 1.690 ;
        RECT  2.610 1.450 2.700 1.670 ;
        RECT  1.770 0.710 1.890 1.800 ;
        RECT  0.130 0.590 0.250 1.880 ;
        RECT  0.870 1.480 1.020 1.640 ;
        RECT  3.340 0.480 3.500 1.910 ;
    END
END MUX3D0

MACRO MUX3D1
    CLASS CORE ;
    FOREIGN MUX3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.960 4.550 2.100 ;
        RECT  4.550 0.420 4.710 2.100 ;
        RECT  4.710 1.960 4.740 2.100 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.490 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.990 0.560 1.515 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.725 0.880 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.520 0.300 ;
        RECT  0.520 -0.300 0.740 0.600 ;
        RECT  0.740 -0.300 2.210 0.300 ;
        RECT  2.210 -0.300 2.430 0.340 ;
        RECT  2.430 -0.300 4.120 0.300 ;
        RECT  4.120 -0.300 4.340 0.340 ;
        RECT  4.340 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 1.970 0.710 2.820 ;
        RECT  0.710 2.220 2.210 2.820 ;
        RECT  2.210 2.180 2.430 2.820 ;
        RECT  2.430 2.220 4.120 2.820 ;
        RECT  4.120 2.180 4.340 2.820 ;
        RECT  4.340 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 1.820 3.970 1.980 ;
        RECT  3.810 0.710 3.970 0.870 ;
        RECT  1.530 0.470 3.000 0.590 ;
        RECT  3.000 0.470 3.160 2.030 ;
        RECT  2.810 1.140 2.880 1.360 ;
        RECT  1.800 0.710 1.890 2.060 ;
        RECT  1.890 1.640 2.020 2.060 ;
        RECT  1.890 0.710 2.040 0.870 ;
        RECT  0.280 0.540 0.360 0.700 ;
        RECT  0.280 1.730 0.910 1.850 ;
        RECT  0.910 1.730 1.030 2.050 ;
        RECT  1.030 1.910 1.460 2.050 ;
        RECT  1.460 1.910 1.680 2.070 ;
        RECT  1.000 0.590 1.150 1.610 ;
        RECT  4.270 0.470 4.430 1.290 ;
        RECT  3.540 0.470 4.270 0.590 ;
        RECT  3.380 0.470 3.540 2.030 ;
        RECT  3.690 0.710 3.810 1.980 ;
        RECT  1.370 0.470 1.530 1.760 ;
        RECT  2.650 0.710 2.810 1.760 ;
        RECT  1.770 0.710 1.800 1.760 ;
        RECT  0.120 0.540 0.280 1.850 ;
        RECT  0.860 1.450 1.000 1.610 ;
    END
END MUX3D1

MACRO MUX3D2
    CLASS CORE ;
    FOREIGN MUX3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.960 4.510 2.100 ;
        RECT  4.510 1.390 4.570 2.100 ;
        RECT  4.510 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.670 2.100 ;
        RECT  4.670 1.960 4.700 2.100 ;
        RECT  4.670 0.780 4.710 1.515 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.490 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.990 0.560 1.515 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 0.725 0.880 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.520 0.300 ;
        RECT  0.520 -0.300 0.740 0.600 ;
        RECT  0.740 -0.300 2.210 0.300 ;
        RECT  2.210 -0.300 2.430 0.340 ;
        RECT  2.430 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 1.970 0.710 2.820 ;
        RECT  0.710 2.220 2.210 2.820 ;
        RECT  2.210 2.180 2.430 2.820 ;
        RECT  2.430 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.280 1.730 0.910 1.850 ;
        RECT  0.910 1.730 1.030 2.050 ;
        RECT  1.030 1.910 1.460 2.050 ;
        RECT  1.460 1.910 1.680 2.100 ;
        RECT  1.000 0.590 1.150 1.610 ;
        RECT  0.280 0.540 0.360 0.700 ;
        RECT  1.890 0.710 2.040 0.870 ;
        RECT  1.890 1.640 2.020 2.060 ;
        RECT  1.800 0.710 1.890 2.060 ;
        RECT  2.810 1.140 2.880 1.360 ;
        RECT  3.000 0.470 3.160 2.030 ;
        RECT  1.530 0.470 3.000 0.590 ;
        RECT  3.810 0.710 3.970 0.870 ;
        RECT  3.810 1.820 3.970 1.980 ;
        RECT  4.350 1.080 4.450 1.240 ;
        RECT  4.230 0.470 4.350 1.240 ;
        RECT  3.540 0.470 4.230 0.590 ;
        RECT  3.380 0.470 3.540 2.030 ;
        RECT  3.690 0.710 3.810 1.980 ;
        RECT  1.370 0.470 1.530 1.760 ;
        RECT  2.650 0.710 2.810 1.760 ;
        RECT  1.770 0.710 1.800 1.760 ;
        RECT  0.120 0.540 0.280 1.850 ;
        RECT  0.860 1.450 1.000 1.610 ;
    END
END MUX3D2

MACRO MUX3D4
    CLASS CORE ;
    FOREIGN MUX3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.000 1.650 6.350 2.030 ;
        RECT  6.000 0.490 6.350 0.870 ;
        RECT  6.350 0.490 6.770 2.030 ;
        RECT  6.770 1.650 6.920 2.030 ;
        RECT  6.770 0.490 6.920 0.870 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.005 3.440 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.005 2.480 1.515 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.350 1.235 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.005 3.110 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.560 0.300 ;
        RECT  0.560 -0.300 0.780 0.340 ;
        RECT  0.780 -0.300 5.610 0.300 ;
        RECT  5.610 -0.300 5.830 0.340 ;
        RECT  5.830 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 5.610 2.820 ;
        RECT  5.610 2.180 5.830 2.820 ;
        RECT  5.830 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.970 0.430 1.190 0.850 ;
        RECT  1.060 1.960 1.090 2.100 ;
        RECT  0.900 1.390 1.060 2.100 ;
        RECT  0.360 0.690 0.970 0.850 ;
        RECT  0.260 1.390 0.900 1.510 ;
        RECT  0.870 1.960 0.900 2.100 ;
        RECT  0.260 0.430 0.360 0.850 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.140 0.430 0.260 2.100 ;
        RECT  0.100 1.390 0.140 2.100 ;
        RECT  2.200 0.710 2.320 0.870 ;
        RECT  2.160 1.650 2.280 1.810 ;
        RECT  2.160 0.710 2.200 1.280 ;
        RECT  2.080 0.710 2.160 1.810 ;
        RECT  2.040 1.120 2.080 1.810 ;
        RECT  2.820 0.710 3.020 0.870 ;
        RECT  2.820 1.890 3.000 2.050 ;
        RECT  2.700 0.710 2.820 2.050 ;
        RECT  1.860 1.930 2.700 2.050 ;
        RECT  1.810 0.710 1.960 0.870 ;
        RECT  1.810 1.410 1.860 2.050 ;
        RECT  1.700 0.710 1.810 2.050 ;
        RECT  3.600 0.710 3.740 1.800 ;
        RECT  3.450 0.710 3.600 0.870 ;
        RECT  3.860 0.470 4.000 2.050 ;
        RECT  1.570 0.470 3.860 0.590 ;
        RECT  1.480 0.470 1.570 0.630 ;
        RECT  4.690 0.710 5.460 0.870 ;
        RECT  5.410 1.960 5.440 2.100 ;
        RECT  5.250 1.390 5.410 2.100 ;
        RECT  4.790 1.390 5.250 1.510 ;
        RECT  5.220 1.960 5.250 2.100 ;
        RECT  4.690 1.390 4.790 2.000 ;
        RECT  5.830 1.070 6.110 1.230 ;
        RECT  5.710 0.470 5.830 1.230 ;
        RECT  4.380 0.470 5.710 0.590 ;
        RECT  4.570 0.710 4.690 2.000 ;
        RECT  1.320 0.470 1.480 1.910 ;
        RECT  4.220 0.470 4.380 2.050 ;
        RECT  3.440 1.640 3.600 1.800 ;
        RECT  1.690 0.710 1.700 1.530 ;
        RECT  1.930 1.120 2.040 1.280 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  6.000 0.490 6.135 0.870 ;
        RECT  6.000 1.650 6.135 2.030 ;
    END
END MUX3D4

MACRO MUX3ND0
    CLASS CORE ;
    FOREIGN MUX3ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.710 3.430 1.980 ;
        RECT  3.430 1.820 3.570 1.980 ;
        RECT  3.430 0.710 3.570 0.870 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.590 1.240 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.015 0.410 1.235 ;
        RECT  0.410 0.725 0.550 1.235 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.180 1.270 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 0.890 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.550 0.300 ;
        RECT  0.550 -0.300 0.770 0.600 ;
        RECT  0.770 -0.300 2.210 0.300 ;
        RECT  2.210 -0.300 2.430 0.340 ;
        RECT  2.430 -0.300 4.130 0.300 ;
        RECT  4.130 -0.300 4.350 0.340 ;
        RECT  4.350 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.960 0.680 2.820 ;
        RECT  0.680 2.220 2.200 2.820 ;
        RECT  2.200 2.180 2.420 2.820 ;
        RECT  2.420 2.220 4.130 2.820 ;
        RECT  4.130 2.180 4.350 2.820 ;
        RECT  4.350 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.010 0.605 1.150 1.600 ;
        RECT  1.540 1.910 1.780 2.070 ;
        RECT  0.920 1.910 1.540 2.050 ;
        RECT  0.800 1.720 0.920 2.050 ;
        RECT  0.260 1.720 0.800 1.840 ;
        RECT  0.230 0.510 0.290 0.730 ;
        RECT  0.230 1.520 0.260 1.840 ;
        RECT  1.880 0.710 1.960 0.850 ;
        RECT  2.840 1.140 2.880 1.360 ;
        RECT  2.720 0.710 2.840 1.710 ;
        RECT  2.600 0.710 2.720 0.870 ;
        RECT  3.000 0.470 3.160 2.030 ;
        RECT  1.530 0.470 3.000 0.590 ;
        RECT  1.370 0.470 1.530 1.760 ;
        RECT  3.810 0.710 3.970 0.870 ;
        RECT  3.810 1.820 3.970 1.980 ;
        RECT  3.690 0.710 3.810 1.980 ;
        RECT  1.270 1.600 1.370 1.760 ;
        RECT  2.600 1.550 2.720 1.710 ;
        RECT  1.720 0.710 1.880 1.760 ;
        RECT  0.100 0.510 0.230 1.840 ;
        RECT  0.830 1.460 1.010 1.600 ;
    END
END MUX3ND0

MACRO MUX3ND1
    CLASS CORE ;
    FOREIGN MUX3ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.160 1.960 5.190 2.100 ;
        RECT  5.190 0.420 5.350 2.100 ;
        RECT  5.350 1.960 5.380 2.100 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.590 1.240 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.015 0.410 1.235 ;
        RECT  0.410 0.725 0.550 1.235 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.285 4.390 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.180 1.270 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 0.890 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.550 0.300 ;
        RECT  0.550 -0.300 0.770 0.600 ;
        RECT  0.770 -0.300 2.210 0.300 ;
        RECT  2.210 -0.300 2.430 0.340 ;
        RECT  2.430 -0.300 4.770 0.300 ;
        RECT  4.770 -0.300 4.990 0.340 ;
        RECT  4.990 -0.300 5.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.960 0.680 2.820 ;
        RECT  0.680 2.220 2.200 2.820 ;
        RECT  2.200 2.180 2.420 2.820 ;
        RECT  2.420 2.220 4.770 2.820 ;
        RECT  4.770 2.180 4.990 2.820 ;
        RECT  4.990 2.220 5.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.550 0.940 4.710 1.290 ;
        RECT  3.810 1.820 3.970 1.980 ;
        RECT  3.810 0.710 3.970 0.870 ;
        RECT  1.370 0.470 1.530 1.760 ;
        RECT  1.530 0.470 3.000 0.590 ;
        RECT  3.000 0.470 3.160 2.030 ;
        RECT  2.600 0.710 2.720 0.870 ;
        RECT  2.720 0.710 2.840 1.710 ;
        RECT  2.840 1.140 2.880 1.360 ;
        RECT  1.890 0.710 1.970 0.850 ;
        RECT  0.230 1.520 0.260 1.840 ;
        RECT  0.230 0.510 0.290 0.730 ;
        RECT  0.260 1.720 0.800 1.840 ;
        RECT  0.800 1.720 0.920 2.050 ;
        RECT  0.920 1.910 1.540 2.050 ;
        RECT  1.540 1.910 1.780 2.070 ;
        RECT  1.010 0.605 1.150 1.600 ;
        RECT  4.220 0.940 4.550 1.060 ;
        RECT  4.100 0.470 4.220 1.060 ;
        RECT  3.540 0.470 4.100 0.590 ;
        RECT  4.910 0.660 5.070 1.760 ;
        RECT  4.350 0.660 4.910 0.820 ;
        RECT  4.590 1.640 4.910 1.760 ;
        RECT  3.380 0.470 3.540 2.030 ;
        RECT  3.690 0.710 3.810 1.980 ;
        RECT  1.270 1.600 1.370 1.760 ;
        RECT  2.600 1.550 2.720 1.710 ;
        RECT  1.730 0.710 1.890 1.760 ;
        RECT  0.100 0.510 0.230 1.840 ;
        RECT  0.830 1.460 1.010 1.600 ;
        RECT  4.370 1.640 4.590 2.090 ;
    END
END MUX3ND1

MACRO MUX3ND2
    CLASS CORE ;
    FOREIGN MUX3ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.090 1.960 5.120 2.100 ;
        RECT  5.120 1.390 5.210 2.100 ;
        RECT  5.120 0.420 5.210 0.900 ;
        RECT  5.210 0.420 5.280 2.100 ;
        RECT  5.280 1.960 5.310 2.100 ;
        RECT  5.280 0.780 5.350 1.515 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.590 1.240 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.015 0.410 1.235 ;
        RECT  0.410 0.725 0.550 1.235 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.285 4.390 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.180 1.270 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 0.890 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.550 0.300 ;
        RECT  0.550 -0.300 0.770 0.600 ;
        RECT  0.770 -0.300 2.210 0.300 ;
        RECT  2.210 -0.300 2.430 0.340 ;
        RECT  2.430 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.960 0.680 2.820 ;
        RECT  0.680 2.220 2.200 2.820 ;
        RECT  2.200 2.180 2.420 2.820 ;
        RECT  2.420 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.720 0.710 2.840 1.710 ;
        RECT  2.840 1.140 2.880 1.360 ;
        RECT  1.880 0.710 1.960 0.850 ;
        RECT  0.230 1.520 0.260 1.840 ;
        RECT  0.230 0.510 0.290 0.730 ;
        RECT  0.260 1.720 0.800 1.840 ;
        RECT  0.800 1.720 0.920 2.050 ;
        RECT  0.920 1.910 1.540 2.050 ;
        RECT  1.540 1.910 1.780 2.070 ;
        RECT  1.010 0.605 1.150 1.600 ;
        RECT  2.600 0.710 2.720 0.870 ;
        RECT  3.000 0.470 3.160 2.030 ;
        RECT  1.530 0.470 3.000 0.590 ;
        RECT  1.370 0.470 1.530 1.760 ;
        RECT  3.810 0.710 3.970 0.870 ;
        RECT  3.810 1.820 3.970 1.980 ;
        RECT  4.530 0.975 4.690 1.290 ;
        RECT  4.220 0.975 4.530 1.095 ;
        RECT  4.100 0.470 4.220 1.095 ;
        RECT  3.540 0.470 4.100 0.590 ;
        RECT  4.930 1.050 5.030 1.270 ;
        RECT  4.810 0.660 4.930 1.760 ;
        RECT  4.350 0.660 4.810 0.820 ;
        RECT  4.590 1.640 4.810 1.760 ;
        RECT  4.370 1.640 4.590 2.090 ;
        RECT  3.380 0.470 3.540 2.030 ;
        RECT  3.690 0.710 3.810 1.980 ;
        RECT  1.270 1.600 1.370 1.760 ;
        RECT  2.600 1.550 2.720 1.710 ;
        RECT  1.720 0.710 1.880 1.760 ;
        RECT  0.100 0.510 0.230 1.840 ;
        RECT  0.830 1.460 1.010 1.600 ;
    END
END MUX3ND2

MACRO MUX3ND4
    CLASS CORE ;
    FOREIGN MUX3ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.880 1.650 7.310 2.030 ;
        RECT  6.880 0.490 7.310 0.870 ;
        RECT  7.310 0.490 7.730 2.030 ;
        RECT  7.730 1.650 7.840 2.030 ;
        RECT  7.730 0.490 7.840 0.870 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.750 1.515 ;
        RECT  3.750 1.050 3.880 1.270 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END S0
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.800 ;
        RECT  0.690 -0.300 1.270 0.300 ;
        RECT  1.270 -0.300 1.490 0.520 ;
        RECT  1.490 -0.300 3.520 0.300 ;
        RECT  3.520 -0.300 3.740 0.340 ;
        RECT  3.740 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.000 0.690 2.820 ;
        RECT  0.690 2.220 1.270 2.820 ;
        RECT  1.270 2.000 1.490 2.820 ;
        RECT  1.490 2.220 2.740 2.820 ;
        RECT  2.740 2.180 2.960 2.820 ;
        RECT  2.960 2.220 3.520 2.820 ;
        RECT  3.520 2.180 3.740 2.820 ;
        RECT  3.740 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.730 0.640 1.850 1.640 ;
        RECT  0.850 0.640 1.730 0.800 ;
        RECT  2.260 1.930 2.500 2.090 ;
        RECT  1.805 1.930 2.260 2.050 ;
        RECT  1.685 1.760 1.805 2.050 ;
        RECT  0.260 1.760 1.685 1.880 ;
        RECT  2.800 0.710 3.370 0.870 ;
        RECT  3.320 1.960 3.350 2.100 ;
        RECT  3.160 1.390 3.320 2.100 ;
        RECT  2.800 1.390 3.160 1.510 ;
        RECT  3.130 1.960 3.160 2.100 ;
        RECT  2.680 0.710 2.800 1.710 ;
        RECT  2.470 0.710 2.680 0.860 ;
        RECT  4.140 1.080 4.220 1.300 ;
        RECT  4.020 0.710 4.140 1.660 ;
        RECT  3.900 0.710 4.020 0.870 ;
        RECT  4.340 0.470 4.460 2.030 ;
        RECT  4.300 0.470 4.340 0.900 ;
        RECT  4.300 1.790 4.340 2.030 ;
        RECT  2.200 0.470 4.300 0.590 ;
        RECT  6.070 1.030 6.230 1.480 ;
        RECT  4.840 1.360 6.070 1.480 ;
        RECT  6.350 0.750 6.470 1.720 ;
        RECT  6.000 0.750 6.350 0.870 ;
        RECT  6.000 1.600 6.350 1.720 ;
        RECT  5.780 0.450 6.000 0.870 ;
        RECT  5.780 1.600 6.000 2.050 ;
        RECT  5.010 0.710 5.780 0.870 ;
        RECT  5.220 1.600 5.780 1.720 ;
        RECT  6.710 1.080 6.990 1.240 ;
        RECT  6.590 0.470 6.710 2.000 ;
        RECT  6.120 0.470 6.590 0.630 ;
        RECT  6.120 1.840 6.590 2.000 ;
        RECT  5.060 1.600 5.220 2.030 ;
        RECT  4.680 0.660 4.840 2.030 ;
        RECT  2.040 0.470 2.200 1.800 ;
        RECT  3.900 1.500 4.020 1.660 ;
        RECT  2.370 1.550 2.680 1.710 ;
        RECT  0.100 0.590 0.260 1.880 ;
        RECT  0.850 1.480 1.730 1.640 ;
        LAYER M1 ;
        RECT  6.880 0.490 7.095 0.870 ;
        RECT  6.880 1.650 7.095 2.030 ;
    END
END MUX3ND4

MACRO MUX4D0
    CLASS CORE ;
    FOREIGN MUX4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.470 0.660 6.630 2.100 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.005 6.000 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.080 4.250 1.240 ;
        RECT  4.250 1.005 4.390 1.515 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.590 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 4.090 0.300 ;
        RECT  4.090 -0.300 4.310 0.340 ;
        RECT  4.310 -0.300 6.020 0.300 ;
        RECT  6.020 -0.300 6.240 0.340 ;
        RECT  6.240 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 2.570 2.820 ;
        RECT  2.570 2.180 2.790 2.820 ;
        RECT  2.790 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 6.020 2.820 ;
        RECT  6.020 2.180 6.240 2.820 ;
        RECT  6.240 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.420 0.470 6.190 0.590 ;
        RECT  6.190 0.470 6.350 1.290 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  5.600 0.710 5.720 2.030 ;
        RECT  5.720 1.640 5.870 1.800 ;
        RECT  5.720 0.710 5.880 0.870 ;
        RECT  3.310 0.760 3.440 0.920 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  4.880 1.495 4.920 1.735 ;
        RECT  4.880 0.470 4.920 0.790 ;
        RECT  4.920 0.470 5.040 1.735 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  3.810 0.760 4.030 0.900 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.760 3.070 0.920 ;
        RECT  3.070 0.760 3.190 1.570 ;
        RECT  1.890 0.760 1.990 0.920 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  5.260 0.470 5.420 1.735 ;
        RECT  1.390 0.710 1.550 1.810 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  4.520 0.710 4.680 1.665 ;
        RECT  3.690 0.760 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.760 1.890 1.570 ;
        RECT  0.870 1.635 1.030 1.795 ;
    END
END MUX4D0

MACRO MUX4D1
    CLASS CORE ;
    FOREIGN MUX4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.440 1.960 6.470 2.100 ;
        RECT  6.470 0.420 6.630 2.100 ;
        RECT  6.630 1.960 6.660 2.100 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.005 6.000 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.530 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 6.020 0.300 ;
        RECT  6.020 -0.300 6.240 0.340 ;
        RECT  6.240 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 6.020 2.820 ;
        RECT  6.020 2.180 6.240 2.820 ;
        RECT  6.240 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.420 0.470 6.190 0.590 ;
        RECT  6.190 0.470 6.350 1.290 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  5.600 0.710 5.720 2.030 ;
        RECT  5.720 1.640 5.850 1.800 ;
        RECT  5.720 0.710 5.880 0.870 ;
        RECT  3.310 0.740 3.440 0.900 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  4.880 1.570 4.920 1.790 ;
        RECT  4.880 0.470 4.920 0.740 ;
        RECT  4.920 0.470 5.040 1.790 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  3.810 0.740 4.030 0.880 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.740 3.070 0.900 ;
        RECT  3.070 0.740 3.190 1.570 ;
        RECT  1.890 0.740 1.990 0.900 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  1.390 0.710 1.550 1.810 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  4.520 0.710 4.680 1.730 ;
        RECT  3.690 0.740 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.740 1.890 1.570 ;
        RECT  0.750 1.635 1.030 1.795 ;
        RECT  5.260 0.470 5.420 1.790 ;
    END
END MUX4D1

MACRO MUX4D2
    CLASS CORE ;
    FOREIGN MUX4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.350 1.960 6.380 2.100 ;
        RECT  6.380 1.390 6.470 2.100 ;
        RECT  6.380 0.420 6.470 0.900 ;
        RECT  6.470 0.420 6.540 2.100 ;
        RECT  6.540 1.960 6.570 2.100 ;
        RECT  6.540 0.725 6.630 1.515 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.005 6.000 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.530 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  5.600 0.710 5.720 2.030 ;
        RECT  5.720 1.640 5.850 1.800 ;
        RECT  5.720 0.710 5.880 0.870 ;
        RECT  3.310 0.740 3.440 0.900 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  4.880 1.570 4.920 1.790 ;
        RECT  4.880 0.470 4.920 0.740 ;
        RECT  4.920 0.470 5.040 1.790 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  3.810 0.740 4.030 0.880 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.740 3.070 0.900 ;
        RECT  3.070 0.740 3.190 1.570 ;
        RECT  1.890 0.740 1.990 0.900 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  6.240 1.050 6.320 1.270 ;
        RECT  6.130 0.735 6.240 1.270 ;
        RECT  6.120 0.470 6.130 1.270 ;
        RECT  6.010 0.470 6.120 0.855 ;
        RECT  5.420 0.470 6.010 0.590 ;
        RECT  5.260 0.470 5.420 1.790 ;
        RECT  1.390 0.710 1.550 1.810 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  4.520 0.710 4.680 1.730 ;
        RECT  3.690 0.740 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.740 1.890 1.570 ;
        RECT  0.750 1.635 1.030 1.795 ;
    END
END MUX4D2

MACRO MUX4D4
    CLASS CORE ;
    FOREIGN MUX4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.060 1.650 9.550 2.030 ;
        RECT  9.060 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 2.030 ;
        RECT  9.970 1.650 10.070 2.030 ;
        RECT  9.970 0.490 10.070 0.870 ;
        END
    END Z
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 6.950 1.515 ;
        RECT  6.950 1.050 7.100 1.270 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.630 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.610 ;
        RECT  0.670 -0.300 3.670 0.300 ;
        RECT  3.670 -0.300 3.890 0.640 ;
        RECT  3.890 -0.300 9.450 0.300 ;
        RECT  9.450 -0.300 9.670 0.340 ;
        RECT  9.670 -0.300 10.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.220 2.820 ;
        RECT  1.220 2.180 1.440 2.820 ;
        RECT  1.440 2.220 2.880 2.820 ;
        RECT  2.880 2.180 3.100 2.820 ;
        RECT  3.100 2.220 3.710 2.820 ;
        RECT  3.710 2.180 3.930 2.820 ;
        RECT  3.930 2.220 4.530 2.820 ;
        RECT  4.530 2.180 4.750 2.820 ;
        RECT  4.750 2.220 6.020 2.820 ;
        RECT  6.020 2.180 6.240 2.820 ;
        RECT  6.240 2.220 6.800 2.820 ;
        RECT  6.800 2.180 7.020 2.820 ;
        RECT  7.020 2.220 9.450 2.820 ;
        RECT  9.450 2.180 9.670 2.820 ;
        RECT  9.670 2.220 10.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.050 0.720 5.170 1.570 ;
        RECT  2.550 0.720 3.310 0.880 ;
        RECT  2.550 1.430 3.530 1.570 ;
        RECT  0.810 1.640 1.600 1.800 ;
        RECT  1.170 0.810 1.600 0.930 ;
        RECT  1.600 0.810 1.640 1.800 ;
        RECT  1.640 0.710 1.760 1.800 ;
        RECT  1.760 0.710 1.880 0.870 ;
        RECT  4.250 0.720 5.050 0.880 ;
        RECT  5.040 1.930 5.280 2.090 ;
        RECT  2.490 1.930 5.040 2.050 ;
        RECT  5.040 0.430 5.280 0.590 ;
        RECT  4.130 0.470 5.040 0.590 ;
        RECT  4.010 0.470 4.130 0.880 ;
        RECT  3.550 0.760 4.010 0.880 ;
        RECT  3.430 0.470 3.550 0.880 ;
        RECT  2.400 0.470 3.430 0.590 ;
        RECT  2.180 0.430 2.400 0.590 ;
        RECT  0.910 0.470 2.180 0.590 ;
        RECT  1.700 1.930 1.940 2.090 ;
        RECT  0.530 1.930 1.700 2.050 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  5.790 0.710 6.700 0.870 ;
        RECT  6.440 1.430 6.600 1.670 ;
        RECT  5.790 1.430 6.440 1.570 ;
        RECT  7.380 1.050 7.500 1.270 ;
        RECT  7.620 0.470 7.740 1.810 ;
        RECT  7.580 0.470 7.620 0.740 ;
        RECT  7.580 1.570 7.620 1.810 ;
        RECT  5.540 0.470 7.580 0.590 ;
        RECT  5.420 0.470 5.540 1.570 ;
        RECT  5.290 0.740 5.420 0.900 ;
        RECT  8.420 0.710 8.580 0.870 ;
        RECT  8.420 1.640 8.550 1.800 ;
        RECT  8.300 0.710 8.420 2.050 ;
        RECT  5.630 1.930 8.300 2.050 ;
        RECT  5.510 1.690 5.630 2.050 ;
        RECT  2.210 1.690 5.510 1.810 ;
        RECT  8.940 1.080 9.335 1.240 ;
        RECT  8.820 0.470 8.940 1.240 ;
        RECT  8.120 0.470 8.820 0.590 ;
        RECT  2.050 0.710 2.210 1.810 ;
        RECT  5.290 1.430 5.420 1.570 ;
        RECT  7.220 0.710 7.380 1.730 ;
        RECT  5.670 0.710 5.790 1.570 ;
        RECT  7.960 0.470 8.120 1.810 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.250 1.930 2.490 2.090 ;
        RECT  4.100 1.430 5.050 1.570 ;
        RECT  2.430 0.720 2.550 1.570 ;
        RECT  1.030 0.710 1.170 0.930 ;
        LAYER M1 ;
        RECT  9.060 1.650 9.335 2.030 ;
        RECT  9.060 0.490 9.335 0.870 ;
    END
END MUX4D4

MACRO MUX4ND0
    CLASS CORE ;
    FOREIGN MUX4ND0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.570 5.350 1.715 ;
        RECT  5.350 1.495 5.420 1.715 ;
        RECT  5.350 0.570 5.420 0.790 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.005 6.000 1.515 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.080 4.250 1.240 ;
        RECT  4.250 1.005 4.390 1.515 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.590 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 4.090 0.300 ;
        RECT  4.090 -0.300 4.310 0.340 ;
        RECT  4.310 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 2.570 2.820 ;
        RECT  2.570 2.180 2.790 2.820 ;
        RECT  2.790 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  5.600 0.710 5.720 2.030 ;
        RECT  5.720 1.640 5.870 1.800 ;
        RECT  5.720 0.710 5.880 0.870 ;
        RECT  3.310 0.760 3.440 0.920 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  4.880 1.495 4.920 1.735 ;
        RECT  4.880 0.470 4.920 0.790 ;
        RECT  4.920 0.470 5.040 1.735 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  3.810 0.760 4.030 0.920 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.870 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.760 3.070 0.920 ;
        RECT  3.070 0.760 3.190 1.570 ;
        RECT  1.890 0.760 1.990 0.920 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  4.520 0.710 4.680 1.665 ;
        RECT  3.690 0.760 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.760 1.890 1.570 ;
        RECT  0.870 1.635 1.030 1.795 ;
        RECT  1.390 0.710 1.550 1.810 ;
    END
END MUX4ND0

MACRO MUX4ND1
    CLASS CORE ;
    FOREIGN MUX4ND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.960 6.790 2.100 ;
        RECT  6.790 0.420 6.950 2.100 ;
        RECT  6.950 1.960 6.980 2.100 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.910 6.060 2.070 ;
        RECT  6.060 1.910 6.490 2.050 ;
        RECT  6.490 1.565 6.630 2.075 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.530 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.000 0.470 6.230 0.630 ;
        RECT  6.230 0.470 6.350 1.760 ;
        RECT  6.350 1.050 6.670 1.270 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  5.600 1.585 5.710 2.030 ;
        RECT  5.710 1.380 5.720 2.030 ;
        RECT  5.720 1.380 5.830 1.745 ;
        RECT  5.620 0.710 5.860 0.870 ;
        RECT  5.830 1.380 5.990 1.500 ;
        RECT  5.860 0.750 5.990 0.870 ;
        RECT  5.990 0.750 6.110 1.500 ;
        RECT  5.420 1.040 5.870 1.260 ;
        RECT  3.310 0.740 3.440 0.900 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  4.880 1.570 4.920 1.790 ;
        RECT  4.880 0.470 4.920 0.740 ;
        RECT  4.920 0.470 5.040 1.790 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  3.810 0.740 4.030 0.880 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.740 3.070 0.900 ;
        RECT  3.070 0.740 3.190 1.570 ;
        RECT  1.890 0.740 1.990 0.900 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  6.000 1.620 6.230 1.760 ;
        RECT  1.390 0.710 1.550 1.810 ;
        RECT  5.260 0.500 5.420 1.790 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  4.520 0.710 4.680 1.730 ;
        RECT  3.690 0.740 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.740 1.890 1.570 ;
        RECT  0.750 1.635 1.030 1.795 ;
    END
END MUX4ND1

MACRO MUX4ND2
    CLASS CORE ;
    FOREIGN MUX4ND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.760 1.960 6.790 2.100 ;
        RECT  6.790 0.420 6.950 2.100 ;
        RECT  6.950 1.960 6.980 2.100 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.840 1.910 6.060 2.070 ;
        RECT  6.060 1.910 6.490 2.050 ;
        RECT  6.490 1.565 6.630 2.075 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.530 ;
        RECT  0.670 -0.300 2.350 0.300 ;
        RECT  2.350 -0.300 2.570 0.640 ;
        RECT  2.570 -0.300 7.160 0.300 ;
        RECT  7.160 -0.300 7.410 0.340 ;
        RECT  7.410 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.160 2.820 ;
        RECT  2.160 2.180 2.380 2.820 ;
        RECT  2.380 2.220 4.090 2.820 ;
        RECT  4.090 2.180 4.310 2.820 ;
        RECT  4.310 2.220 7.160 2.820 ;
        RECT  7.160 2.180 7.410 2.820 ;
        RECT  7.410 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 0.740 4.030 0.880 ;
        RECT  1.700 1.930 3.180 2.050 ;
        RECT  3.180 1.930 3.400 2.090 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 1.930 1.140 2.050 ;
        RECT  1.140 1.930 1.360 2.090 ;
        RECT  0.910 0.470 1.520 0.590 ;
        RECT  1.520 0.430 1.740 0.590 ;
        RECT  1.740 0.470 2.110 0.590 ;
        RECT  2.110 0.470 2.230 0.880 ;
        RECT  2.230 0.760 2.690 0.880 ;
        RECT  2.690 0.470 2.810 0.880 ;
        RECT  2.810 0.470 3.060 0.590 ;
        RECT  3.060 0.430 3.300 0.590 ;
        RECT  2.930 0.740 3.070 0.900 ;
        RECT  3.070 0.740 3.190 1.570 ;
        RECT  1.890 0.740 1.990 0.900 ;
        RECT  1.890 1.430 2.010 1.570 ;
        RECT  1.030 0.710 1.170 1.795 ;
        RECT  3.810 1.430 3.930 1.570 ;
        RECT  4.680 1.050 4.770 1.270 ;
        RECT  4.920 0.470 5.040 1.790 ;
        RECT  4.880 0.470 4.920 0.740 ;
        RECT  4.880 1.570 4.920 1.790 ;
        RECT  3.560 0.470 4.880 0.590 ;
        RECT  3.440 0.470 3.560 1.570 ;
        RECT  3.310 0.740 3.440 0.900 ;
        RECT  5.420 1.040 5.870 1.260 ;
        RECT  5.990 0.750 6.110 1.500 ;
        RECT  5.860 0.750 5.990 0.870 ;
        RECT  5.830 1.380 5.990 1.500 ;
        RECT  5.620 0.710 5.860 0.870 ;
        RECT  5.720 1.380 5.830 1.745 ;
        RECT  5.710 1.380 5.720 2.030 ;
        RECT  5.600 1.585 5.710 2.030 ;
        RECT  3.650 1.910 5.600 2.030 ;
        RECT  3.530 1.690 3.650 2.030 ;
        RECT  1.550 1.690 3.530 1.810 ;
        RECT  6.350 1.050 6.670 1.270 ;
        RECT  6.230 0.470 6.350 1.760 ;
        RECT  6.000 0.470 6.230 0.630 ;
        RECT  1.390 0.710 1.550 1.810 ;
        RECT  5.260 0.500 5.420 1.790 ;
        RECT  3.310 1.430 3.440 1.570 ;
        RECT  4.520 0.710 4.680 1.730 ;
        RECT  3.690 0.740 3.810 1.570 ;
        RECT  1.480 1.930 1.700 2.090 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.930 1.430 3.070 1.570 ;
        RECT  1.770 0.740 1.890 1.570 ;
        RECT  6.000 1.620 6.230 1.760 ;
        RECT  0.750 1.635 1.030 1.795 ;
    END
END MUX4ND2

MACRO MUX4ND4
    CLASS CORE ;
    FOREIGN MUX4ND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.780 1.650 10.190 2.030 ;
        RECT  9.780 0.490 10.190 0.870 ;
        RECT  10.190 0.490 10.610 2.030 ;
        RECT  10.610 1.650 10.740 2.030 ;
        RECT  10.610 0.490 10.740 0.870 ;
        END
    END ZN
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 6.950 1.515 ;
        RECT  6.950 1.050 7.100 1.270 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END S0
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.630 1.235 ;
        END
    END I3
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END I1
    PIN I0
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.610 ;
        RECT  0.670 -0.300 3.670 0.300 ;
        RECT  3.670 -0.300 3.890 0.640 ;
        RECT  3.890 -0.300 9.380 0.300 ;
        RECT  9.380 -0.300 9.600 0.340 ;
        RECT  9.600 -0.300 11.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.220 2.820 ;
        RECT  1.220 2.180 1.440 2.820 ;
        RECT  1.440 2.220 2.880 2.820 ;
        RECT  2.880 2.180 3.100 2.820 ;
        RECT  3.100 2.220 3.710 2.820 ;
        RECT  3.710 2.180 3.930 2.820 ;
        RECT  3.930 2.220 4.530 2.820 ;
        RECT  4.530 2.180 4.750 2.820 ;
        RECT  4.750 2.220 6.020 2.820 ;
        RECT  6.020 2.180 6.240 2.820 ;
        RECT  6.240 2.220 6.800 2.820 ;
        RECT  6.800 2.180 7.020 2.820 ;
        RECT  7.020 2.220 9.380 2.820 ;
        RECT  9.380 2.180 9.600 2.820 ;
        RECT  9.600 2.220 11.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.010 0.470 4.130 0.880 ;
        RECT  4.130 0.470 5.040 0.590 ;
        RECT  5.040 0.430 5.280 0.590 ;
        RECT  2.490 1.930 5.040 2.050 ;
        RECT  5.040 1.930 5.280 2.090 ;
        RECT  4.250 0.720 5.050 0.880 ;
        RECT  5.050 0.720 5.170 1.570 ;
        RECT  2.550 0.720 3.310 0.880 ;
        RECT  2.550 1.430 3.530 1.570 ;
        RECT  0.810 1.640 1.600 1.800 ;
        RECT  1.170 0.810 1.600 0.930 ;
        RECT  1.600 0.810 1.640 1.800 ;
        RECT  1.640 0.710 1.760 1.800 ;
        RECT  1.760 0.710 1.880 0.870 ;
        RECT  3.550 0.760 4.010 0.880 ;
        RECT  3.430 0.470 3.550 0.880 ;
        RECT  2.400 0.470 3.430 0.590 ;
        RECT  2.180 0.430 2.400 0.590 ;
        RECT  0.910 0.470 2.180 0.590 ;
        RECT  1.700 1.930 1.940 2.090 ;
        RECT  0.530 1.930 1.700 2.050 ;
        RECT  0.790 0.470 0.910 0.850 ;
        RECT  0.530 0.730 0.790 0.850 ;
        RECT  0.410 0.730 0.530 2.050 ;
        RECT  0.330 0.730 0.410 0.850 ;
        RECT  0.070 1.890 0.410 2.050 ;
        RECT  0.210 0.420 0.330 0.850 ;
        RECT  5.790 0.710 6.700 0.870 ;
        RECT  6.440 1.430 6.600 1.670 ;
        RECT  5.790 1.430 6.440 1.570 ;
        RECT  7.380 1.050 7.500 1.270 ;
        RECT  7.620 0.470 7.740 1.810 ;
        RECT  7.580 0.470 7.620 0.740 ;
        RECT  7.580 1.570 7.620 1.810 ;
        RECT  5.540 0.470 7.580 0.590 ;
        RECT  5.420 0.470 5.540 1.570 ;
        RECT  5.290 0.740 5.420 0.900 ;
        RECT  8.120 1.080 9.150 1.240 ;
        RECT  9.300 0.750 9.420 1.480 ;
        RECT  8.500 0.750 9.300 0.870 ;
        RECT  8.500 1.360 9.300 1.480 ;
        RECT  8.340 0.500 8.500 0.870 ;
        RECT  8.340 1.360 8.500 2.050 ;
        RECT  5.630 1.930 8.340 2.050 ;
        RECT  5.510 1.690 5.630 2.050 ;
        RECT  2.210 1.690 5.510 1.810 ;
        RECT  9.660 1.080 9.880 1.240 ;
        RECT  9.540 0.470 9.660 1.760 ;
        RECT  8.970 0.470 9.540 0.630 ;
        RECT  9.210 1.600 9.540 1.760 ;
        RECT  2.050 0.710 2.210 1.810 ;
        RECT  7.960 0.500 8.120 1.810 ;
        RECT  5.290 1.430 5.420 1.570 ;
        RECT  7.220 0.710 7.380 1.730 ;
        RECT  5.670 0.710 5.790 1.570 ;
        RECT  8.990 1.600 9.210 2.020 ;
        RECT  0.070 0.420 0.210 0.580 ;
        RECT  2.250 1.930 2.490 2.090 ;
        RECT  4.100 1.430 5.050 1.570 ;
        RECT  2.430 0.720 2.550 1.570 ;
        RECT  1.030 0.710 1.170 0.930 ;
        LAYER M1 ;
        RECT  9.780 1.650 9.975 2.030 ;
        RECT  9.780 0.490 9.975 0.870 ;
    END
END MUX4ND4

MACRO ND2D0
    CLASS CORE ;
    FOREIGN ND2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.710 0.560 1.720 ;
        RECT  0.560 0.710 0.890 0.870 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.610 2.820 ;
        RECT  0.610 2.180 0.830 2.820 ;
        RECT  0.830 2.220 0.960 2.820 ;
        END
    END VDD
END ND2D0

MACRO ND2D1
    CLASS CORE ;
    FOREIGN ND2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.960 0.400 2.100 ;
        RECT  0.400 0.715 0.560 2.100 ;
        RECT  0.560 1.960 0.590 2.100 ;
        RECT  0.560 0.715 0.670 0.840 ;
        RECT  0.670 0.420 0.890 0.840 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.960 2.820 ;
        END
    END VDD
END ND2D1

MACRO ND2D2
    CLASS CORE ;
    FOREIGN ND2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.665 0.550 1.760 ;
        RECT  0.550 0.665 1.090 0.825 ;
        RECT  0.550 1.600 1.440 1.760 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 2.030 ;
        RECT  0.250 1.890 1.560 2.030 ;
        RECT  1.330 1.080 1.560 1.240 ;
        RECT  1.560 1.080 1.680 2.030 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.190 0.300 ;
        RECT  0.190 -0.300 0.410 0.340 ;
        RECT  0.410 -0.300 1.510 0.300 ;
        RECT  1.510 -0.300 1.730 0.340 ;
        RECT  1.730 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
END ND2D2

MACRO ND2D3
    CLASS CORE ;
    FOREIGN ND2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.440 0.470 0.560 1.810 ;
        RECT  0.560 1.410 0.660 1.810 ;
        RECT  0.660 1.410 1.130 1.540 ;
        RECT  1.130 1.410 1.350 1.810 ;
        RECT  1.870 1.425 2.290 1.935 ;
        RECT  2.290 1.425 2.330 1.550 ;
        RECT  0.560 0.470 2.330 0.630 ;
        RECT  2.330 0.470 2.470 1.550 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 2.050 ;
        RECT  0.250 1.930 1.470 2.050 ;
        RECT  1.470 1.030 1.630 2.050 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.070 1.235 ;
        RECT  1.070 0.750 1.190 1.235 ;
        RECT  1.190 0.750 2.050 0.870 ;
        RECT  2.050 0.750 2.210 1.230 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.170 0.300 ;
        RECT  0.170 -0.300 0.390 0.340 ;
        RECT  0.390 -0.300 1.500 0.300 ;
        RECT  1.500 -0.300 1.720 0.340 ;
        RECT  1.720 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.520 2.820 ;
        RECT  1.520 2.180 1.740 2.820 ;
        RECT  1.740 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.440 0.470 0.560 1.810 ;
        RECT  0.560 1.410 0.660 1.810 ;
        RECT  0.660 1.410 1.130 1.540 ;
        RECT  1.130 1.410 1.350 1.810 ;
        RECT  0.560 0.470 2.330 0.630 ;
        RECT  2.330 0.470 2.470 1.210 ;
    END
END ND2D3

MACRO ND2D4
    CLASS CORE ;
    FOREIGN ND2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.710 0.550 2.040 ;
        RECT  0.550 0.710 1.050 0.870 ;
        RECT  0.550 1.880 2.510 2.040 ;
        RECT  2.140 0.710 2.510 0.870 ;
        RECT  2.510 0.710 2.630 2.040 ;
        RECT  2.630 1.425 2.930 2.040 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.470 0.250 1.290 ;
        RECT  0.250 0.470 1.520 0.590 ;
        RECT  1.520 0.470 1.680 1.290 ;
        RECT  1.680 0.470 2.950 0.590 ;
        RECT  2.950 0.470 3.110 1.255 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.070 1.235 ;
        RECT  1.070 1.005 1.190 1.560 ;
        RECT  1.190 1.440 2.040 1.560 ;
        RECT  2.040 1.030 2.200 1.560 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 1.500 0.300 ;
        RECT  1.500 -0.300 1.720 0.340 ;
        RECT  1.720 -0.300 2.820 0.300 ;
        RECT  2.820 -0.300 3.040 0.340 ;
        RECT  3.040 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.510 0.710 2.630 1.210 ;
        RECT  0.550 1.880 2.295 2.040 ;
        RECT  0.550 0.710 1.050 0.870 ;
        RECT  0.430 0.710 0.550 2.040 ;
        RECT  2.140 0.710 2.510 0.870 ;
    END
END ND2D4

MACRO ND2D8
    CLASS CORE ;
    FOREIGN ND2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.650 0.740 2.030 ;
        RECT  0.740 0.710 0.860 2.030 ;
        RECT  0.860 0.710 1.210 0.870 ;
        RECT  0.860 1.650 2.495 2.030 ;
        RECT  2.280 0.710 2.495 0.870 ;
        RECT  2.495 0.710 2.615 2.030 ;
        RECT  2.615 1.650 2.830 2.030 ;
        RECT  2.830 1.425 3.250 2.030 ;
        RECT  3.250 1.650 3.570 2.030 ;
        RECT  3.570 0.710 3.690 2.030 ;
        RECT  3.690 0.710 3.930 0.870 ;
        RECT  3.690 1.650 5.310 2.030 ;
        RECT  5.000 0.710 5.310 0.870 ;
        RECT  5.310 0.710 5.430 2.030 ;
        RECT  5.430 1.650 5.630 2.030 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.470 0.570 1.290 ;
        RECT  0.570 0.470 1.630 0.590 ;
        RECT  1.630 0.470 1.750 1.240 ;
        RECT  1.750 1.080 1.870 1.240 ;
        RECT  1.750 0.470 2.750 0.590 ;
        RECT  2.750 0.470 2.870 1.180 ;
        RECT  2.870 1.020 3.330 1.180 ;
        RECT  3.330 0.470 3.450 1.180 ;
        RECT  4.350 1.080 4.470 1.240 ;
        RECT  3.450 0.470 4.470 0.590 ;
        RECT  4.470 0.470 4.590 1.240 ;
        RECT  4.590 0.470 5.550 0.590 ;
        RECT  5.550 0.470 5.710 1.290 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.390 1.235 ;
        RECT  1.390 1.005 1.510 1.480 ;
        RECT  1.510 1.360 2.215 1.480 ;
        RECT  2.215 1.030 2.375 1.480 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.310 0.300 ;
        RECT  0.310 -0.300 0.530 0.340 ;
        RECT  0.530 -0.300 1.640 0.300 ;
        RECT  1.640 -0.300 1.860 0.340 ;
        RECT  1.860 -0.300 2.990 0.300 ;
        RECT  2.990 -0.300 3.210 0.750 ;
        RECT  3.210 -0.300 4.350 0.300 ;
        RECT  4.350 -0.300 4.570 0.340 ;
        RECT  4.570 -0.300 5.680 0.300 ;
        RECT  5.680 -0.300 5.900 0.340 ;
        RECT  5.900 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.170 2.820 ;
        RECT  0.170 2.180 0.390 2.820 ;
        RECT  0.390 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.030 1.030 5.190 1.480 ;
        RECT  3.970 1.360 5.030 1.480 ;
        RECT  3.810 1.030 3.970 1.480 ;
        LAYER M1 ;
        RECT  2.280 0.710 2.495 0.870 ;
        RECT  2.495 0.710 2.615 2.030 ;
        RECT  3.570 0.710 3.690 2.030 ;
        RECT  3.690 0.710 3.930 0.870 ;
        RECT  3.690 1.650 5.310 2.030 ;
        RECT  5.000 0.710 5.310 0.870 ;
        RECT  5.310 0.710 5.430 2.030 ;
        RECT  5.430 1.650 5.630 2.030 ;
        RECT  0.860 1.650 2.495 2.030 ;
        RECT  0.860 0.710 1.210 0.870 ;
        RECT  0.740 0.710 0.860 2.030 ;
        RECT  0.580 1.650 0.740 2.030 ;
        RECT  3.465 1.650 3.570 2.030 ;
    END
END ND2D8

MACRO ND3D0
    CLASS CORE ;
    FOREIGN ND3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.500 1.820 1.350 1.980 ;
        RECT  1.150 0.520 1.350 0.680 ;
        RECT  1.350 0.520 1.510 1.980 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.535 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.260 0.300 ;
        RECT  0.260 -0.300 0.480 0.340 ;
        RECT  0.480 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.920 2.820 ;
        RECT  0.920 2.180 1.140 2.820 ;
        RECT  1.140 2.220 1.600 2.820 ;
        END
    END VDD
END ND3D0

MACRO ND3D1
    CLASS CORE ;
    FOREIGN ND3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.640 0.740 2.060 ;
        RECT  0.740 1.640 1.310 1.800 ;
        RECT  1.310 1.640 1.370 2.060 ;
        RECT  1.170 0.430 1.370 0.850 ;
        RECT  1.370 0.430 1.390 2.060 ;
        RECT  1.390 0.730 1.510 2.060 ;
        RECT  1.510 1.640 1.530 2.060 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.190 0.300 ;
        RECT  0.190 -0.300 0.410 0.340 ;
        RECT  0.410 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.920 2.820 ;
        RECT  0.920 2.180 1.140 2.820 ;
        RECT  1.140 2.220 1.600 2.820 ;
        END
    END VDD
END ND3D1

MACRO ND3D2
    CLASS CORE ;
    FOREIGN ND3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.450 1.390 0.870 ;
        RECT  0.430 1.880 2.330 2.040 ;
        RECT  1.390 0.750 2.330 0.870 ;
        RECT  2.330 0.750 2.470 2.040 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.760 ;
        RECT  0.550 1.640 2.015 1.760 ;
        RECT  2.015 1.030 2.175 1.760 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        RECT  0.880 1.395 1.680 1.515 ;
        RECT  1.680 1.030 1.840 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.180 0.300 ;
        RECT  0.180 -0.300 0.400 0.340 ;
        RECT  0.400 -0.300 2.160 0.300 ;
        RECT  2.160 -0.300 2.380 0.340 ;
        RECT  2.380 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.560 2.820 ;
        END
    END VDD
END ND3D2

MACRO ND3D3
    CLASS CORE ;
    FOREIGN ND3D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.120 0.480 0.240 2.040 ;
        RECT  0.240 0.480 1.360 0.640 ;
        RECT  0.240 1.880 2.830 2.040 ;
        RECT  2.830 1.425 3.250 2.040 ;
        RECT  3.250 1.425 3.330 1.585 ;
        RECT  3.230 0.420 3.330 0.900 ;
        RECT  3.330 0.420 3.390 1.585 ;
        RECT  3.390 0.780 3.450 1.585 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.050 0.550 1.760 ;
        RECT  0.550 1.640 2.310 1.760 ;
        RECT  2.310 1.005 2.470 1.760 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.395 1.580 1.515 ;
        RECT  1.580 1.080 1.700 1.515 ;
        RECT  1.700 1.080 1.940 1.240 ;
        RECT  1.940 0.750 2.060 1.240 ;
        RECT  2.060 0.750 2.690 0.870 ;
        RECT  2.690 0.750 2.850 1.250 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.820 1.310 1.270 ;
        RECT  1.310 0.820 1.700 0.940 ;
        RECT  1.700 0.480 1.820 0.940 ;
        RECT  1.820 0.480 2.970 0.600 ;
        RECT  2.970 0.480 3.110 1.230 ;
        RECT  3.110 1.040 3.210 1.200 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 2.140 0.300 ;
        RECT  2.140 -0.300 2.360 0.340 ;
        RECT  2.360 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.420 3.330 0.900 ;
        RECT  0.120 0.480 0.240 2.040 ;
        RECT  0.240 0.480 1.360 0.640 ;
        RECT  0.240 1.880 2.615 2.040 ;
        RECT  3.330 0.420 3.390 1.210 ;
        RECT  3.390 0.780 3.450 1.210 ;
    END
END ND3D3

MACRO ND3D4
    CLASS CORE ;
    FOREIGN ND3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.110 0.470 0.230 1.680 ;
        RECT  0.230 1.560 0.450 1.680 ;
        RECT  0.450 1.560 0.610 2.040 ;
        RECT  0.230 0.470 1.130 0.590 ;
        RECT  1.130 0.430 1.370 0.590 ;
        RECT  3.160 0.430 3.400 0.590 ;
        RECT  0.610 1.880 3.790 2.040 ;
        RECT  3.790 1.425 4.210 2.040 ;
        RECT  4.210 1.425 4.260 1.650 ;
        RECT  3.400 0.470 4.260 0.590 ;
        RECT  4.260 0.470 4.380 1.650 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 0.710 0.510 1.270 ;
        RECT  0.510 0.710 2.000 0.830 ;
        RECT  2.000 0.710 2.160 1.270 ;
        RECT  2.160 0.710 4.000 0.830 ;
        RECT  4.000 0.710 4.140 1.210 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.080 0.740 1.240 ;
        RECT  0.740 0.950 0.860 1.760 ;
        RECT  0.860 0.950 1.630 1.070 ;
        RECT  1.630 0.950 1.790 1.270 ;
        RECT  2.330 1.005 2.710 1.235 ;
        RECT  2.710 0.950 2.830 1.235 ;
        RECT  0.860 1.640 3.440 1.760 ;
        RECT  2.830 0.950 3.440 1.070 ;
        RECT  3.440 0.950 3.560 1.760 ;
        RECT  3.560 1.020 3.870 1.180 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.190 1.270 1.515 ;
        RECT  1.270 1.285 1.510 1.515 ;
        RECT  1.510 1.395 3.100 1.515 ;
        RECT  3.100 1.190 3.220 1.515 ;
        RECT  3.220 1.190 3.320 1.330 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.140 0.300 ;
        RECT  0.140 -0.300 0.360 0.340 ;
        RECT  0.360 -0.300 2.110 0.300 ;
        RECT  2.110 -0.300 2.330 0.340 ;
        RECT  2.330 -0.300 4.130 0.300 ;
        RECT  4.130 -0.300 4.350 0.340 ;
        RECT  4.350 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.270 2.820 ;
        RECT  4.270 2.180 4.490 2.820 ;
        RECT  4.490 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.160 0.430 3.400 0.590 ;
        RECT  0.110 0.470 0.230 1.680 ;
        RECT  0.230 1.560 0.450 1.680 ;
        RECT  0.450 1.560 0.610 2.040 ;
        RECT  0.230 0.470 1.130 0.590 ;
        RECT  1.130 0.430 1.370 0.590 ;
        RECT  0.610 1.880 3.575 2.040 ;
        RECT  3.400 0.470 4.260 0.590 ;
        RECT  4.260 0.470 4.380 1.210 ;
    END
END ND3D4

MACRO ND3D8
    CLASS CORE ;
    FOREIGN ND3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.960 0.480 2.100 ;
        RECT  0.480 1.370 0.640 2.100 ;
        RECT  0.640 1.930 0.670 2.100 ;
        RECT  0.670 1.930 1.170 2.050 ;
        RECT  1.170 1.930 1.200 2.100 ;
        RECT  1.200 1.370 1.360 2.100 ;
        RECT  1.360 1.930 1.390 2.100 ;
        RECT  1.390 1.930 1.900 2.050 ;
        RECT  1.900 1.930 1.930 2.100 ;
        RECT  1.930 1.370 2.090 2.100 ;
        RECT  2.090 1.930 2.120 2.100 ;
        RECT  2.120 1.930 2.630 2.050 ;
        RECT  2.630 1.930 2.660 2.100 ;
        RECT  2.660 1.370 2.820 2.100 ;
        RECT  2.820 1.930 2.850 2.100 ;
        RECT  2.850 1.930 3.410 2.050 ;
        RECT  3.410 1.930 3.440 2.100 ;
        RECT  3.440 1.370 3.600 2.100 ;
        RECT  3.600 1.930 3.630 2.100 ;
        RECT  3.630 1.930 4.190 2.050 ;
        RECT  4.190 1.930 4.220 2.100 ;
        RECT  4.220 1.370 4.380 2.100 ;
        RECT  4.380 1.930 4.410 2.100 ;
        RECT  4.410 1.930 4.970 2.050 ;
        RECT  4.970 1.930 5.000 2.100 ;
        RECT  5.000 1.370 5.160 2.100 ;
        RECT  5.160 1.930 5.190 2.100 ;
        RECT  5.190 1.930 5.750 2.050 ;
        RECT  5.750 1.930 5.780 2.100 ;
        RECT  5.780 1.370 5.940 2.100 ;
        RECT  5.940 1.930 5.970 2.100 ;
        RECT  5.970 1.930 6.530 2.050 ;
        RECT  6.530 1.930 6.560 2.100 ;
        RECT  6.560 1.370 6.720 2.100 ;
        RECT  6.720 1.930 6.750 2.100 ;
        RECT  6.750 1.930 7.310 2.050 ;
        RECT  7.310 1.930 7.340 2.100 ;
        RECT  7.340 1.370 7.500 2.100 ;
        RECT  7.500 1.930 7.530 2.100 ;
        RECT  7.530 1.930 8.090 2.050 ;
        RECT  8.090 1.930 8.120 2.100 ;
        RECT  8.120 1.370 8.280 2.100 ;
        RECT  8.280 1.930 8.310 2.100 ;
        RECT  8.310 1.930 8.590 2.050 ;
        RECT  6.630 0.710 8.590 0.870 ;
        RECT  8.590 0.710 9.010 2.050 ;
        RECT  9.010 1.670 9.090 2.050 ;
        RECT  9.010 0.710 9.170 0.870 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.005 7.910 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 3.800 2.820 ;
        RECT  3.800 2.180 4.020 2.820 ;
        RECT  4.020 2.220 4.580 2.820 ;
        RECT  4.580 2.180 4.800 2.820 ;
        RECT  4.800 2.220 5.360 2.820 ;
        RECT  5.360 2.180 5.580 2.820 ;
        RECT  5.580 2.220 6.140 2.820 ;
        RECT  6.140 2.180 6.360 2.820 ;
        RECT  6.360 2.220 6.920 2.820 ;
        RECT  6.920 2.180 7.140 2.820 ;
        RECT  7.140 2.220 7.700 2.820 ;
        RECT  7.700 2.180 7.920 2.820 ;
        RECT  7.920 2.220 8.480 2.820 ;
        RECT  8.480 2.180 8.700 2.820 ;
        RECT  8.700 2.220 9.260 2.820 ;
        RECT  9.260 2.180 9.480 2.820 ;
        RECT  9.480 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.910 0.720 6.150 0.880 ;
        RECT  5.370 0.760 5.910 0.880 ;
        RECT  5.150 0.720 5.370 0.880 ;
        RECT  4.610 0.760 5.150 0.880 ;
        RECT  4.390 0.720 4.610 0.880 ;
        RECT  3.850 0.760 4.390 0.880 ;
        RECT  3.630 0.720 3.850 0.880 ;
        RECT  3.090 0.760 3.630 0.880 ;
        RECT  2.870 0.450 3.090 0.880 ;
        RECT  2.390 0.760 2.870 0.880 ;
        RECT  2.170 0.450 2.390 0.880 ;
        RECT  1.690 0.760 2.170 0.880 ;
        RECT  1.470 0.450 1.690 0.880 ;
        RECT  0.990 0.760 1.470 0.880 ;
        RECT  0.770 0.450 0.990 0.880 ;
        RECT  0.290 0.760 0.770 0.880 ;
        RECT  9.310 0.470 9.530 0.900 ;
        RECT  8.770 0.470 9.310 0.590 ;
        RECT  8.550 0.430 8.770 0.590 ;
        RECT  8.010 0.470 8.550 0.590 ;
        RECT  7.790 0.430 8.010 0.590 ;
        RECT  7.250 0.470 7.790 0.590 ;
        RECT  7.030 0.430 7.250 0.590 ;
        RECT  6.490 0.470 7.030 0.590 ;
        RECT  6.270 0.470 6.490 0.900 ;
        RECT  5.750 0.470 6.270 0.590 ;
        RECT  5.530 0.430 5.750 0.590 ;
        RECT  4.990 0.470 5.530 0.590 ;
        RECT  4.770 0.430 4.990 0.590 ;
        RECT  4.230 0.470 4.770 0.590 ;
        RECT  4.010 0.430 4.230 0.590 ;
        RECT  3.470 0.470 4.010 0.590 ;
        RECT  3.230 0.430 3.470 0.590 ;
        RECT  0.070 0.450 0.290 0.880 ;
        LAYER M1 ;
        RECT  6.750 1.930 7.310 2.050 ;
        RECT  7.310 1.930 7.340 2.100 ;
        RECT  7.340 1.370 7.500 2.100 ;
        RECT  7.500 1.930 7.530 2.100 ;
        RECT  7.530 1.930 8.090 2.050 ;
        RECT  8.090 1.930 8.120 2.100 ;
        RECT  8.120 1.370 8.280 2.100 ;
        RECT  8.280 1.930 8.310 2.100 ;
        RECT  8.310 1.930 8.375 2.050 ;
        RECT  6.720 1.930 6.750 2.100 ;
        RECT  6.560 1.370 6.720 2.100 ;
        RECT  6.530 1.930 6.560 2.100 ;
        RECT  5.970 1.930 6.530 2.050 ;
        RECT  5.940 1.930 5.970 2.100 ;
        RECT  5.780 1.370 5.940 2.100 ;
        RECT  5.750 1.930 5.780 2.100 ;
        RECT  5.190 1.930 5.750 2.050 ;
        RECT  5.160 1.930 5.190 2.100 ;
        RECT  5.000 1.370 5.160 2.100 ;
        RECT  4.970 1.930 5.000 2.100 ;
        RECT  4.410 1.930 4.970 2.050 ;
        RECT  4.380 1.930 4.410 2.100 ;
        RECT  4.220 1.370 4.380 2.100 ;
        RECT  4.190 1.930 4.220 2.100 ;
        RECT  3.630 1.930 4.190 2.050 ;
        RECT  3.600 1.930 3.630 2.100 ;
        RECT  3.440 1.370 3.600 2.100 ;
        RECT  3.410 1.930 3.440 2.100 ;
        RECT  2.850 1.930 3.410 2.050 ;
        RECT  2.820 1.930 2.850 2.100 ;
        RECT  2.660 1.370 2.820 2.100 ;
        RECT  2.630 1.930 2.660 2.100 ;
        RECT  2.120 1.930 2.630 2.050 ;
        RECT  2.090 1.930 2.120 2.100 ;
        RECT  1.930 1.370 2.090 2.100 ;
        RECT  1.900 1.930 1.930 2.100 ;
        RECT  1.390 1.930 1.900 2.050 ;
        RECT  1.360 1.930 1.390 2.100 ;
        RECT  1.200 1.370 1.360 2.100 ;
        RECT  1.170 1.930 1.200 2.100 ;
        RECT  0.670 1.930 1.170 2.050 ;
        RECT  0.640 1.930 0.670 2.100 ;
        RECT  0.480 1.370 0.640 2.100 ;
        RECT  6.630 0.710 8.375 0.870 ;
        RECT  0.450 1.960 0.480 2.100 ;
    END
END ND3D8

MACRO ND4D0
    CLASS CORE ;
    FOREIGN ND4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.870 1.690 2.030 ;
        RECT  1.470 0.460 1.690 0.620 ;
        RECT  1.690 0.460 1.830 2.030 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.005 1.540 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.200 0.300 ;
        RECT  0.200 -0.300 0.420 0.340 ;
        RECT  0.420 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
END ND4D0

MACRO ND4D1
    CLASS CORE ;
    FOREIGN ND4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.650 0.700 2.070 ;
        RECT  0.700 1.650 1.220 1.770 ;
        RECT  1.220 1.650 1.440 2.070 ;
        RECT  1.440 1.650 1.690 1.770 ;
        RECT  1.490 0.430 1.690 0.850 ;
        RECT  1.690 0.430 1.710 1.770 ;
        RECT  1.710 0.730 1.830 1.770 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.200 0.300 ;
        RECT  0.200 -0.300 0.420 0.340 ;
        RECT  0.420 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.920 2.820 ;
        END
    END VDD
END ND4D1

MACRO ND4D2
    CLASS CORE ;
    FOREIGN ND4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.750 0.550 1.515 ;
        RECT  0.570 1.960 0.600 2.100 ;
        RECT  0.550 1.390 0.600 1.515 ;
        RECT  0.550 0.750 0.710 0.910 ;
        RECT  0.600 1.390 0.760 2.100 ;
        RECT  0.760 1.930 0.790 2.100 ;
        RECT  0.790 1.930 1.400 2.050 ;
        RECT  1.400 1.930 1.430 2.100 ;
        RECT  1.430 1.370 1.590 2.100 ;
        RECT  1.590 1.930 1.620 2.100 ;
        RECT  1.620 1.930 2.230 2.050 ;
        RECT  2.230 1.930 2.260 2.100 ;
        RECT  2.260 1.370 2.420 2.100 ;
        RECT  2.420 1.930 2.450 2.100 ;
        RECT  2.450 1.930 3.060 2.050 ;
        RECT  3.060 1.635 3.280 2.050 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.005 3.440 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.140 0.300 ;
        RECT  3.140 -0.300 3.360 0.340 ;
        RECT  3.360 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.160 2.820 ;
        RECT  0.160 2.180 0.380 2.820 ;
        RECT  0.380 2.220 0.980 2.820 ;
        RECT  0.980 2.180 1.200 2.820 ;
        RECT  1.200 2.220 1.810 2.820 ;
        RECT  1.810 2.180 2.030 2.820 ;
        RECT  2.030 2.220 2.640 2.820 ;
        RECT  2.640 2.180 2.860 2.820 ;
        RECT  2.860 2.220 3.470 2.820 ;
        RECT  3.470 2.180 3.690 2.820 ;
        RECT  3.690 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.610 0.470 1.830 0.630 ;
        RECT  1.070 0.470 1.610 0.590 ;
        RECT  0.850 0.470 1.070 0.885 ;
        RECT  2.350 0.710 2.590 0.870 ;
        RECT  1.450 0.750 2.350 0.870 ;
        RECT  3.550 0.470 3.770 0.890 ;
        RECT  2.950 0.470 3.550 0.590 ;
        RECT  2.730 0.470 2.950 0.890 ;
        RECT  2.190 0.470 2.730 0.590 ;
        RECT  1.970 0.470 2.190 0.630 ;
        RECT  1.210 0.710 1.450 0.870 ;
        RECT  0.070 0.470 0.850 0.630 ;
    END
END ND4D2

MACRO ND4D3
    CLASS CORE ;
    FOREIGN ND4D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.450 0.290 0.880 ;
        RECT  0.070 1.640 0.590 2.020 ;
        RECT  0.290 0.760 0.590 0.880 ;
        RECT  0.590 0.760 1.010 2.020 ;
        RECT  1.010 0.760 1.050 0.880 ;
        RECT  1.010 1.640 5.050 2.020 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.005 4.400 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.910 0.300 ;
        RECT  3.910 -0.300 4.130 0.340 ;
        RECT  4.130 -0.300 4.730 0.300 ;
        RECT  4.730 -0.300 4.950 0.340 ;
        RECT  4.950 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.250 2.820 ;
        RECT  1.250 2.180 1.470 2.820 ;
        RECT  1.470 2.220 2.040 2.820 ;
        RECT  2.040 2.180 2.260 2.820 ;
        RECT  2.260 2.220 2.830 2.820 ;
        RECT  2.830 2.180 3.050 2.820 ;
        RECT  3.050 2.220 3.630 2.820 ;
        RECT  3.630 2.180 3.850 2.820 ;
        RECT  3.850 2.220 4.430 2.820 ;
        RECT  4.430 2.180 4.650 2.820 ;
        RECT  4.650 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.400 0.470 2.210 0.630 ;
        RECT  1.240 0.470 1.400 0.940 ;
        RECT  2.570 0.750 3.350 0.870 ;
        RECT  2.350 0.440 2.570 0.870 ;
        RECT  4.320 0.470 4.540 0.880 ;
        RECT  3.710 0.470 4.320 0.630 ;
        RECT  3.490 0.470 3.710 0.890 ;
        RECT  2.710 0.470 3.490 0.630 ;
        RECT  1.570 0.750 2.350 0.870 ;
        RECT  0.430 0.470 1.240 0.630 ;
        LAYER M1 ;
        RECT  0.290 0.760 0.375 0.880 ;
        RECT  0.070 1.640 0.375 2.020 ;
        RECT  0.070 0.450 0.290 0.880 ;
        RECT  1.225 1.640 5.050 2.020 ;
    END
END ND4D3

MACRO ND4D4
    CLASS CORE ;
    FOREIGN ND4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.650 0.910 2.030 ;
        RECT  0.510 0.760 0.910 0.920 ;
        RECT  0.910 0.760 1.330 2.030 ;
        RECT  1.330 1.650 1.510 2.030 ;
        RECT  1.330 0.760 1.530 0.920 ;
        RECT  1.510 1.880 2.050 2.030 ;
        RECT  2.050 1.635 2.270 2.030 ;
        RECT  2.270 1.880 2.810 2.030 ;
        RECT  2.810 1.620 3.030 2.030 ;
        RECT  3.030 1.880 3.910 2.030 ;
        RECT  3.910 1.620 4.130 2.030 ;
        RECT  4.130 1.880 4.670 2.030 ;
        RECT  4.670 1.620 4.890 2.030 ;
        RECT  4.890 1.880 5.360 2.030 ;
        RECT  5.360 1.635 5.580 2.030 ;
        RECT  5.580 1.880 6.050 2.030 ;
        RECT  6.050 1.620 6.270 2.030 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.520 1.005 5.680 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.240 1.005 4.400 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.000 1.005 2.160 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        RECT  0.230 1.080 0.505 1.240 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.370 0.470 3.410 0.590 ;
        RECT  6.430 0.470 6.650 0.890 ;
        RECT  5.960 0.470 6.430 0.630 ;
        RECT  5.740 0.470 5.960 0.890 ;
        RECT  5.270 0.470 5.740 0.630 ;
        RECT  5.050 0.470 5.270 0.890 ;
        RECT  3.530 0.470 5.050 0.630 ;
        RECT  2.030 0.750 4.910 0.885 ;
        RECT  0.150 0.470 0.370 0.880 ;
        LAYER M1 ;
        RECT  6.050 1.620 6.270 2.030 ;
        RECT  5.580 1.880 6.050 2.030 ;
        RECT  5.360 1.635 5.580 2.030 ;
        RECT  4.890 1.880 5.360 2.030 ;
        RECT  4.670 1.620 4.890 2.030 ;
        RECT  4.130 1.880 4.670 2.030 ;
        RECT  3.910 1.620 4.130 2.030 ;
        RECT  3.030 1.880 3.910 2.030 ;
        RECT  2.810 1.620 3.030 2.030 ;
        RECT  2.270 1.880 2.810 2.030 ;
        RECT  2.050 1.635 2.270 2.030 ;
        RECT  0.510 0.760 0.695 0.920 ;
        RECT  0.530 1.650 0.695 2.030 ;
        RECT  1.545 1.880 2.050 2.030 ;
    END
END ND4D4

MACRO ND4D8
    CLASS CORE ;
    FOREIGN ND4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.640 2.830 2.020 ;
        RECT  1.920 0.760 2.830 0.900 ;
        RECT  2.830 0.760 3.250 2.020 ;
        RECT  3.250 1.640 4.260 2.020 ;
        RECT  3.250 0.760 4.280 0.900 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.565 1.150 1.795 ;
        RECT  1.150 1.030 1.310 1.795 ;
        RECT  1.310 1.565 1.510 1.795 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.285 0.810 1.795 ;
        RECT  0.810 1.030 0.870 1.795 ;
        RECT  0.870 1.030 0.970 1.405 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.080 1.005 0.240 1.515 ;
        END
    END A1
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.510 1.050 1.690 1.270 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END A4
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.145 2.820 ;
        RECT  0.145 2.180 0.365 2.820 ;
        RECT  0.365 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.640 1.050 4.700 1.270 ;
        RECT  4.520 0.470 4.640 1.270 ;
        RECT  1.690 0.470 4.520 0.590 ;
        RECT  1.570 0.470 1.690 0.870 ;
        RECT  0.535 0.750 1.570 0.870 ;
        RECT  1.250 1.930 1.490 2.090 ;
        RECT  0.780 1.930 1.250 2.050 ;
        RECT  0.535 1.930 0.780 2.070 ;
        RECT  0.530 0.750 0.535 2.070 ;
        RECT  0.415 0.450 0.530 2.070 ;
        RECT  5.610 1.960 5.640 2.100 ;
        RECT  5.450 0.420 5.610 0.900 ;
        RECT  5.450 1.390 5.610 2.100 ;
        RECT  4.940 0.780 5.450 0.900 ;
        RECT  4.940 1.390 5.450 1.510 ;
        RECT  5.420 1.960 5.450 2.100 ;
        RECT  4.920 1.960 4.950 2.100 ;
        RECT  4.920 0.780 4.940 1.510 ;
        RECT  4.820 0.420 4.920 2.100 ;
        RECT  4.760 0.420 4.820 0.900 ;
        RECT  4.760 1.390 4.820 2.100 ;
        RECT  4.320 1.390 4.760 1.510 ;
        RECT  4.730 1.960 4.760 2.100 ;
        RECT  4.160 1.030 4.320 1.510 ;
        RECT  0.310 0.450 0.415 0.880 ;
        LAYER M1 ;
        RECT  1.920 0.760 2.615 0.900 ;
        RECT  1.940 1.640 2.615 2.020 ;
        RECT  3.465 0.760 4.280 0.900 ;
        RECT  3.465 1.640 4.260 2.020 ;
    END
END ND4D8

MACRO NR2D0
    CLASS CORE ;
    FOREIGN NR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.660 0.560 1.800 ;
        RECT  0.560 1.640 0.900 1.800 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.610 0.300 ;
        RECT  0.610 -0.300 0.830 0.340 ;
        RECT  0.830 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 0.960 2.820 ;
        END
    END VDD
END NR2D0

MACRO NR2D1
    CLASS CORE ;
    FOREIGN NR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 0.420 0.560 1.760 ;
        RECT  0.560 1.640 0.680 1.760 ;
        RECT  0.680 1.640 0.900 2.060 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.960 2.820 ;
        END
    END VDD
END NR2D1

MACRO NR2D2
    CLASS CORE ;
    FOREIGN NR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 0.460 0.690 0.880 ;
        RECT  0.830 1.640 1.050 1.800 ;
        RECT  0.690 0.720 1.050 0.880 ;
        RECT  1.050 0.720 1.190 1.800 ;
        RECT  1.190 0.720 1.230 0.880 ;
        RECT  1.230 0.460 1.450 0.880 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 2.040 ;
        RECT  0.560 1.920 1.360 2.040 ;
        RECT  1.360 1.030 1.520 2.040 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.190 2.820 ;
        RECT  0.190 2.180 0.410 2.820 ;
        RECT  0.410 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 1.920 2.820 ;
        END
    END VDD
END NR2D2

MACRO NR2D3
    CLASS CORE ;
    FOREIGN NR2D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 0.450 0.670 0.610 ;
        RECT  0.670 0.470 0.720 0.610 ;
        RECT  0.720 0.470 0.840 1.550 ;
        RECT  0.840 0.470 0.860 1.810 ;
        RECT  0.860 1.410 1.060 1.810 ;
        RECT  0.860 0.470 1.170 0.600 ;
        RECT  1.170 0.450 1.390 0.600 ;
        RECT  1.390 0.470 1.920 0.600 ;
        RECT  1.920 0.450 2.140 0.600 ;
        RECT  1.870 1.425 2.290 1.935 ;
        RECT  2.290 1.425 2.370 1.585 ;
        RECT  2.140 0.470 2.370 0.600 ;
        RECT  2.370 0.470 2.490 1.585 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 2.050 ;
        RECT  0.550 1.930 1.360 2.050 ;
        RECT  1.360 1.030 1.520 2.050 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 0.725 1.190 1.290 ;
        RECT  1.190 0.725 2.030 0.845 ;
        RECT  2.030 0.725 2.250 1.180 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.430 0.450 0.670 0.610 ;
        RECT  0.670 0.470 0.720 0.610 ;
        RECT  0.720 0.470 0.840 1.550 ;
        RECT  0.840 0.470 0.860 1.810 ;
        RECT  0.860 1.410 1.060 1.810 ;
        RECT  0.860 0.470 1.170 0.600 ;
        RECT  1.170 0.450 1.390 0.600 ;
        RECT  1.390 0.470 1.920 0.600 ;
        RECT  1.920 0.450 2.140 0.600 ;
        RECT  2.140 0.470 2.370 0.600 ;
        RECT  2.370 0.470 2.490 1.210 ;
    END
END NR2D3

MACRO NR2D4
    CLASS CORE ;
    FOREIGN NR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.710 0.550 1.790 ;
        RECT  0.550 1.630 0.810 1.790 ;
        RECT  0.810 1.630 1.030 2.050 ;
        RECT  0.550 0.710 1.360 0.870 ;
        RECT  1.030 1.630 2.510 1.790 ;
        RECT  2.510 1.425 2.630 1.935 ;
        RECT  1.810 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.770 1.935 ;
        RECT  2.770 1.425 2.930 1.935 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.470 0.250 1.290 ;
        RECT  0.250 0.470 1.520 0.590 ;
        RECT  1.520 0.470 1.680 1.270 ;
        RECT  1.680 0.470 2.950 0.590 ;
        RECT  2.950 0.470 3.110 1.255 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.070 1.235 ;
        RECT  1.070 1.005 1.190 1.510 ;
        RECT  1.190 1.390 2.040 1.510 ;
        RECT  2.040 1.030 2.200 1.510 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.480 2.820 ;
        RECT  1.480 2.180 1.700 2.820 ;
        RECT  1.700 2.220 2.800 2.820 ;
        RECT  2.800 2.180 3.020 2.820 ;
        RECT  3.020 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.630 0.710 2.770 1.210 ;
        RECT  1.030 1.630 2.295 1.790 ;
        RECT  0.550 0.710 1.360 0.870 ;
        RECT  0.810 1.630 1.030 2.050 ;
        RECT  0.550 1.630 0.810 1.790 ;
        RECT  0.410 0.710 0.550 1.790 ;
        RECT  1.810 0.710 2.630 0.870 ;
    END
END NR2D4

MACRO NR2D8
    CLASS CORE ;
    FOREIGN NR2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.380 3.670 1.810 ;
        RECT  3.670 1.380 4.210 1.500 ;
        RECT  4.210 1.380 4.430 1.810 ;
        RECT  0.470 0.500 4.430 0.880 ;
        RECT  4.430 0.500 4.850 1.500 ;
        RECT  4.850 1.380 4.970 1.500 ;
        RECT  4.970 1.380 5.190 1.810 ;
        RECT  5.190 1.380 5.730 1.500 ;
        RECT  4.850 0.500 5.920 0.880 ;
        RECT  5.730 1.380 5.950 1.810 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.150 1.005 6.310 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.110 1.640 6.330 2.050 ;
        RECT  5.570 1.930 6.110 2.050 ;
        RECT  5.350 1.620 5.570 2.050 ;
        RECT  4.810 1.930 5.350 2.050 ;
        RECT  4.590 1.620 4.810 2.050 ;
        RECT  4.050 1.930 4.590 2.050 ;
        RECT  3.830 1.620 4.050 2.050 ;
        RECT  3.290 1.930 3.830 2.050 ;
        RECT  3.260 1.930 3.290 2.100 ;
        RECT  3.100 1.370 3.260 2.100 ;
        RECT  3.070 1.930 3.100 2.100 ;
        RECT  2.540 1.930 3.070 2.050 ;
        RECT  2.510 1.930 2.540 2.100 ;
        RECT  2.350 1.370 2.510 2.100 ;
        RECT  2.320 1.930 2.350 2.100 ;
        RECT  1.790 1.930 2.320 2.050 ;
        RECT  1.760 1.930 1.790 2.100 ;
        RECT  1.600 1.370 1.760 2.100 ;
        RECT  1.570 1.930 1.600 2.100 ;
        RECT  1.040 1.930 1.570 2.050 ;
        RECT  1.010 1.930 1.040 2.100 ;
        RECT  0.850 1.370 1.010 2.100 ;
        RECT  0.820 1.930 0.850 2.100 ;
        RECT  0.290 1.930 0.820 2.050 ;
        RECT  0.260 1.930 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  5.730 1.380 5.950 1.810 ;
        RECT  5.190 1.380 5.730 1.500 ;
        RECT  3.670 1.380 4.210 1.500 ;
        RECT  0.470 0.500 4.215 0.880 ;
        RECT  3.450 1.380 3.670 1.810 ;
        RECT  5.065 0.500 5.920 0.880 ;
        RECT  5.065 1.380 5.190 1.810 ;
    END
END NR2D8

MACRO NR3D0
    CLASS CORE ;
    FOREIGN NR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.490 0.470 1.340 0.630 ;
        RECT  1.150 1.640 1.370 2.060 ;
        RECT  1.340 0.470 1.370 0.690 ;
        RECT  1.370 0.470 1.510 1.760 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.220 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.120 0.300 ;
        RECT  0.120 -0.300 0.340 0.340 ;
        RECT  0.340 -0.300 0.910 0.300 ;
        RECT  0.910 -0.300 1.130 0.340 ;
        RECT  1.130 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 1.600 2.820 ;
        END
    END VDD
END NR3D0

MACRO NR3D1
    CLASS CORE ;
    FOREIGN NR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.710 0.550 1.810 ;
        RECT  0.550 1.650 1.100 1.810 ;
        RECT  1.100 1.650 1.320 2.070 ;
        RECT  0.550 0.710 1.360 0.870 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.470 0.250 1.290 ;
        RECT  0.250 0.470 1.850 0.590 ;
        RECT  1.850 0.430 2.090 0.590 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.030 0.820 1.530 ;
        RECT  0.820 1.410 1.690 1.530 ;
        RECT  1.480 0.710 1.690 0.870 ;
        RECT  1.690 0.710 1.830 1.530 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 2.240 2.820 ;
        END
    END VDD
END NR3D1

MACRO NR3D2
    CLASS CORE ;
    FOREIGN NR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.370 3.430 1.790 ;
        RECT  3.430 1.370 3.790 1.510 ;
        RECT  0.840 0.470 3.790 0.630 ;
        RECT  3.790 0.470 3.970 1.510 ;
        RECT  3.970 0.470 4.190 2.050 ;
        RECT  4.190 0.470 4.210 1.510 ;
        RECT  4.210 0.470 4.420 0.630 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.350 1.235 ;
        RECT  1.350 0.830 1.510 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.310 1.235 ;
        RECT  2.310 0.830 2.470 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.270 1.235 ;
        RECT  3.270 0.830 3.430 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 1.280 0.300 ;
        RECT  1.280 -0.300 1.500 0.340 ;
        RECT  1.500 -0.300 2.110 0.300 ;
        RECT  2.110 -0.300 2.330 0.340 ;
        RECT  2.330 -0.300 2.940 0.300 ;
        RECT  2.940 -0.300 3.160 0.340 ;
        RECT  3.160 -0.300 3.760 0.300 ;
        RECT  3.760 -0.300 3.980 0.340 ;
        RECT  3.980 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.450 1.630 2.670 2.050 ;
        RECT  1.910 1.930 2.450 2.050 ;
        RECT  1.690 1.370 1.910 2.050 ;
        RECT  1.180 1.930 1.690 2.050 ;
        RECT  3.590 1.630 3.810 2.050 ;
        RECT  3.050 1.930 3.590 2.050 ;
        RECT  2.830 1.370 3.050 2.050 ;
        RECT  2.290 1.370 2.830 1.490 ;
        RECT  2.070 1.370 2.290 1.790 ;
        RECT  0.960 1.370 1.180 2.050 ;
        LAYER M1 ;
        RECT  3.430 1.370 3.575 1.510 ;
        RECT  0.840 0.470 3.575 0.630 ;
        RECT  3.210 1.370 3.430 1.790 ;
    END
END NR3D2

MACRO NR3D3
    CLASS CORE ;
    FOREIGN NR3D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.690 1.370 4.750 1.790 ;
        RECT  0.140 0.470 4.750 0.630 ;
        RECT  4.750 0.470 4.910 1.790 ;
        RECT  4.910 0.470 5.170 1.510 ;
        RECT  5.170 1.370 5.450 1.510 ;
        RECT  5.450 1.370 5.670 1.790 ;
        RECT  5.670 1.370 6.210 1.510 ;
        RECT  5.170 0.470 6.210 0.630 ;
        RECT  6.210 1.370 6.430 2.050 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.350 1.235 ;
        RECT  1.350 0.830 1.510 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.005 3.270 1.235 ;
        RECT  3.270 0.830 3.430 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.830 1.235 ;
        RECT  5.830 0.830 5.990 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.580 0.300 ;
        RECT  0.580 -0.300 0.800 0.340 ;
        RECT  0.800 -0.300 1.410 0.300 ;
        RECT  1.410 -0.300 1.630 0.340 ;
        RECT  1.630 -0.300 2.240 0.300 ;
        RECT  2.240 -0.300 2.460 0.340 ;
        RECT  2.460 -0.300 3.070 0.300 ;
        RECT  3.070 -0.300 3.290 0.340 ;
        RECT  3.290 -0.300 3.900 0.300 ;
        RECT  3.900 -0.300 4.120 0.340 ;
        RECT  4.120 -0.300 4.730 0.300 ;
        RECT  4.730 -0.300 4.950 0.340 ;
        RECT  4.950 -0.300 5.550 0.300 ;
        RECT  5.550 -0.300 5.770 0.340 ;
        RECT  5.770 -0.300 6.380 0.300 ;
        RECT  6.380 -0.300 6.600 0.340 ;
        RECT  6.600 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.930 1.630 4.150 2.050 ;
        RECT  3.390 1.930 3.930 2.050 ;
        RECT  3.170 1.630 3.390 2.050 ;
        RECT  2.630 1.930 3.170 2.050 ;
        RECT  2.410 1.370 2.630 2.050 ;
        RECT  1.900 1.930 2.410 2.050 ;
        RECT  1.680 1.370 1.900 2.050 ;
        RECT  1.170 1.930 1.680 2.050 ;
        RECT  5.830 1.630 6.050 2.050 ;
        RECT  5.290 1.930 5.830 2.050 ;
        RECT  5.070 1.630 5.290 2.050 ;
        RECT  4.530 1.930 5.070 2.050 ;
        RECT  4.310 1.370 4.530 2.050 ;
        RECT  3.770 1.370 4.310 1.510 ;
        RECT  3.550 1.370 3.770 1.790 ;
        RECT  3.010 1.370 3.550 1.510 ;
        RECT  2.790 1.370 3.010 1.790 ;
        RECT  0.950 1.370 1.170 2.050 ;
        LAYER M1 ;
        RECT  5.450 1.370 5.670 1.790 ;
        RECT  5.670 1.370 6.210 1.510 ;
        RECT  6.210 1.370 6.430 2.050 ;
        RECT  0.140 0.470 4.535 0.630 ;
        RECT  5.385 0.470 6.210 0.630 ;
        RECT  5.385 1.370 5.450 1.510 ;
    END
END NR3D3

MACRO NR3D4
    CLASS CORE ;
    FOREIGN NR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.900 1.370 6.030 1.790 ;
        RECT  0.760 0.470 6.030 0.630 ;
        RECT  6.030 0.470 6.120 1.790 ;
        RECT  6.120 0.470 6.450 1.490 ;
        RECT  6.450 1.370 6.660 1.490 ;
        RECT  6.660 1.370 6.880 1.790 ;
        RECT  6.880 1.370 7.420 1.490 ;
        RECT  7.420 1.370 7.640 1.790 ;
        RECT  6.450 0.470 7.660 0.630 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.990 1.235 ;
        RECT  1.990 0.830 2.150 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.230 1.235 ;
        RECT  4.230 0.830 4.390 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 7.110 1.235 ;
        RECT  7.110 0.830 7.270 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.370 0.300 ;
        RECT  0.370 -0.300 0.590 0.340 ;
        RECT  0.590 -0.300 1.200 0.300 ;
        RECT  1.200 -0.300 1.420 0.340 ;
        RECT  1.420 -0.300 2.030 0.300 ;
        RECT  2.030 -0.300 2.250 0.340 ;
        RECT  2.250 -0.300 2.860 0.300 ;
        RECT  2.860 -0.300 3.080 0.340 ;
        RECT  3.080 -0.300 3.690 0.300 ;
        RECT  3.690 -0.300 3.910 0.340 ;
        RECT  3.910 -0.300 4.520 0.300 ;
        RECT  4.520 -0.300 4.740 0.340 ;
        RECT  4.740 -0.300 5.350 0.300 ;
        RECT  5.350 -0.300 5.570 0.340 ;
        RECT  5.570 -0.300 6.170 0.300 ;
        RECT  6.170 -0.300 6.390 0.340 ;
        RECT  6.390 -0.300 7.000 0.300 ;
        RECT  7.000 -0.300 7.220 0.340 ;
        RECT  7.220 -0.300 7.830 0.300 ;
        RECT  7.830 -0.300 8.050 0.340 ;
        RECT  8.050 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.170 1.630 5.390 2.050 ;
        RECT  4.630 1.930 5.170 2.050 ;
        RECT  4.410 1.630 4.630 2.050 ;
        RECT  3.870 1.930 4.410 2.050 ;
        RECT  3.650 1.630 3.870 2.050 ;
        RECT  3.110 1.930 3.650 2.050 ;
        RECT  2.890 1.370 3.110 2.050 ;
        RECT  2.350 1.930 2.890 2.050 ;
        RECT  2.130 1.370 2.350 2.050 ;
        RECT  1.590 1.930 2.130 2.050 ;
        RECT  1.370 1.370 1.590 2.050 ;
        RECT  0.830 1.930 1.370 2.050 ;
        RECT  7.800 1.370 8.020 2.050 ;
        RECT  7.260 1.930 7.800 2.050 ;
        RECT  7.040 1.630 7.260 2.050 ;
        RECT  6.500 1.930 7.040 2.050 ;
        RECT  6.280 1.630 6.500 2.050 ;
        RECT  5.740 1.930 6.280 2.050 ;
        RECT  5.520 1.370 5.740 2.050 ;
        RECT  5.010 1.370 5.520 1.490 ;
        RECT  4.790 1.370 5.010 1.790 ;
        RECT  4.250 1.370 4.790 1.490 ;
        RECT  4.030 1.370 4.250 1.790 ;
        RECT  3.490 1.370 4.030 1.490 ;
        RECT  0.610 1.370 0.830 2.050 ;
        RECT  3.270 1.370 3.490 1.790 ;
        LAYER M1 ;
        RECT  7.420 1.370 7.640 1.790 ;
        RECT  6.880 1.370 7.420 1.490 ;
        RECT  0.760 0.470 5.815 0.630 ;
        RECT  6.665 0.470 7.660 0.630 ;
        RECT  6.665 1.370 6.880 1.790 ;
    END
END NR3D4

MACRO NR3D8
    CLASS CORE ;
    FOREIGN NR3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.340 1.370 10.560 1.790 ;
        RECT  10.560 1.370 10.830 1.490 ;
        RECT  0.540 0.470 10.830 0.630 ;
        RECT  10.830 0.470 11.100 1.490 ;
        RECT  11.100 0.470 11.250 1.790 ;
        RECT  11.250 1.370 11.320 1.790 ;
        RECT  11.320 1.370 11.860 1.490 ;
        RECT  11.860 1.370 12.080 1.790 ;
        RECT  12.080 1.370 12.620 1.490 ;
        RECT  12.620 1.370 12.840 1.790 ;
        RECT  12.840 1.370 13.380 1.490 ;
        RECT  13.380 1.370 13.600 1.790 ;
        RECT  13.600 1.370 14.140 1.490 ;
        RECT  14.140 1.370 14.360 1.790 ;
        RECT  11.250 0.470 14.820 0.630 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.630 1.235 ;
        RECT  2.630 0.830 2.790 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.130 1.005 7.430 1.235 ;
        RECT  7.430 0.830 7.590 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  12.250 1.005 12.550 1.235 ;
        RECT  12.550 0.830 12.710 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.150 0.300 ;
        RECT  0.150 -0.300 0.370 0.340 ;
        RECT  0.370 -0.300 0.980 0.300 ;
        RECT  0.980 -0.300 1.200 0.340 ;
        RECT  1.200 -0.300 1.810 0.300 ;
        RECT  1.810 -0.300 2.030 0.340 ;
        RECT  2.030 -0.300 2.640 0.300 ;
        RECT  2.640 -0.300 2.860 0.340 ;
        RECT  2.860 -0.300 3.460 0.300 ;
        RECT  3.460 -0.300 3.680 0.340 ;
        RECT  3.680 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 5.080 0.300 ;
        RECT  5.080 -0.300 5.300 0.340 ;
        RECT  5.300 -0.300 5.880 0.300 ;
        RECT  5.880 -0.300 6.100 0.340 ;
        RECT  6.100 -0.300 6.700 0.300 ;
        RECT  6.700 -0.300 6.920 0.340 ;
        RECT  6.920 -0.300 7.530 0.300 ;
        RECT  7.530 -0.300 7.750 0.340 ;
        RECT  7.750 -0.300 8.360 0.300 ;
        RECT  8.360 -0.300 8.580 0.340 ;
        RECT  8.580 -0.300 9.190 0.300 ;
        RECT  9.190 -0.300 9.410 0.340 ;
        RECT  9.410 -0.300 10.020 0.300 ;
        RECT  10.020 -0.300 10.240 0.340 ;
        RECT  10.240 -0.300 10.850 0.300 ;
        RECT  10.850 -0.300 11.070 0.340 ;
        RECT  11.070 -0.300 11.670 0.300 ;
        RECT  11.670 -0.300 11.890 0.340 ;
        RECT  11.890 -0.300 12.500 0.300 ;
        RECT  12.500 -0.300 12.720 0.340 ;
        RECT  12.720 -0.300 13.330 0.300 ;
        RECT  13.330 -0.300 13.550 0.340 ;
        RECT  13.550 -0.300 14.160 0.300 ;
        RECT  14.160 -0.300 14.380 0.340 ;
        RECT  14.380 -0.300 14.990 0.300 ;
        RECT  14.990 -0.300 15.210 0.340 ;
        RECT  15.210 -0.300 15.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 15.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  9.610 1.630 9.830 2.050 ;
        RECT  9.070 1.930 9.610 2.050 ;
        RECT  8.850 1.630 9.070 2.050 ;
        RECT  8.310 1.930 8.850 2.050 ;
        RECT  8.090 1.630 8.310 2.050 ;
        RECT  7.550 1.930 8.090 2.050 ;
        RECT  7.330 1.630 7.550 2.050 ;
        RECT  6.790 1.930 7.330 2.050 ;
        RECT  6.570 1.630 6.790 2.050 ;
        RECT  6.030 1.930 6.570 2.050 ;
        RECT  5.810 1.630 6.030 2.050 ;
        RECT  5.270 1.930 5.810 2.050 ;
        RECT  5.050 1.370 5.270 2.050 ;
        RECT  4.530 1.930 5.050 2.050 ;
        RECT  4.310 1.370 4.530 2.050 ;
        RECT  3.790 1.930 4.310 2.050 ;
        RECT  3.570 1.370 3.790 2.050 ;
        RECT  3.050 1.930 3.570 2.050 ;
        RECT  2.830 1.370 3.050 2.050 ;
        RECT  2.310 1.930 2.830 2.050 ;
        RECT  2.090 1.370 2.310 2.050 ;
        RECT  1.570 1.930 2.090 2.050 ;
        RECT  1.350 1.370 1.570 2.050 ;
        RECT  0.830 1.930 1.350 2.050 ;
        RECT  14.520 1.370 14.740 2.050 ;
        RECT  13.980 1.930 14.520 2.050 ;
        RECT  13.760 1.630 13.980 2.050 ;
        RECT  13.220 1.930 13.760 2.050 ;
        RECT  13.000 1.630 13.220 2.050 ;
        RECT  12.460 1.930 13.000 2.050 ;
        RECT  12.240 1.630 12.460 2.050 ;
        RECT  11.700 1.930 12.240 2.050 ;
        RECT  11.480 1.630 11.700 2.050 ;
        RECT  10.940 1.930 11.480 2.050 ;
        RECT  10.720 1.630 10.940 2.050 ;
        RECT  10.180 1.930 10.720 2.050 ;
        RECT  9.960 1.370 10.180 2.050 ;
        RECT  9.450 1.370 9.960 1.490 ;
        RECT  9.230 1.370 9.450 1.790 ;
        RECT  8.690 1.370 9.230 1.490 ;
        RECT  8.470 1.370 8.690 1.790 ;
        RECT  7.930 1.370 8.470 1.490 ;
        RECT  7.710 1.370 7.930 1.790 ;
        RECT  7.170 1.370 7.710 1.490 ;
        RECT  6.950 1.370 7.170 1.790 ;
        RECT  6.410 1.370 6.950 1.490 ;
        RECT  6.190 1.370 6.410 1.790 ;
        RECT  5.650 1.370 6.190 1.490 ;
        RECT  5.430 1.370 5.650 1.790 ;
        RECT  0.610 1.370 0.830 2.050 ;
        LAYER M1 ;
        RECT  14.140 1.370 14.360 1.790 ;
        RECT  13.600 1.370 14.140 1.490 ;
        RECT  13.380 1.370 13.600 1.790 ;
        RECT  12.840 1.370 13.380 1.490 ;
        RECT  12.620 1.370 12.840 1.790 ;
        RECT  12.080 1.370 12.620 1.490 ;
        RECT  11.860 1.370 12.080 1.790 ;
        RECT  10.560 1.370 10.615 1.490 ;
        RECT  0.540 0.470 10.615 0.630 ;
        RECT  10.340 1.370 10.560 1.790 ;
        RECT  11.465 0.470 14.820 0.630 ;
        RECT  11.465 1.370 11.860 1.490 ;
    END
END NR3D8

MACRO NR4D0
    CLASS CORE ;
    FOREIGN NR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.640 1.690 2.060 ;
        RECT  0.460 0.470 1.690 0.630 ;
        RECT  1.690 0.470 1.700 2.060 ;
        RECT  1.700 0.470 1.830 1.760 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.190 2.820 ;
        RECT  0.190 2.180 0.410 2.820 ;
        RECT  0.410 2.220 1.920 2.820 ;
        END
    END VDD
END NR4D0

MACRO NR4D1
    CLASS CORE ;
    FOREIGN NR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.410 0.920 1.810 ;
        RECT  0.920 1.410 1.370 1.530 ;
        RECT  0.920 0.660 1.370 0.820 ;
        RECT  1.370 0.660 1.510 1.530 ;
        RECT  1.510 0.660 1.920 0.820 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.560 0.300 ;
        RECT  0.560 -0.300 0.780 0.820 ;
        RECT  0.780 -0.300 2.060 0.300 ;
        RECT  2.060 -0.300 2.280 0.820 ;
        RECT  2.280 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.940 2.820 ;
        RECT  1.940 2.180 2.160 2.820 ;
        RECT  2.160 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.590 1.635 2.810 2.050 ;
        RECT  0.290 1.930 2.590 2.050 ;
        RECT  0.070 1.635 0.290 2.050 ;
    END
END NR4D1

MACRO NR4D2
    CLASS CORE ;
    FOREIGN NR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.480 1.370 4.570 1.790 ;
        RECT  0.450 0.470 4.570 0.630 ;
        RECT  4.570 0.470 4.700 1.790 ;
        RECT  4.700 0.470 4.710 1.490 ;
        RECT  4.710 1.370 5.240 1.490 ;
        RECT  5.240 1.370 5.460 2.050 ;
        RECT  4.710 0.470 5.690 0.630 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 0.830 1.210 1.235 ;
        RECT  1.210 1.005 1.510 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.830 2.490 1.235 ;
        RECT  2.490 1.005 2.790 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 0.830 3.770 1.235 ;
        RECT  3.770 1.005 4.070 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 0.830 5.050 1.235 ;
        RECT  5.050 1.005 5.350 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.890 0.300 ;
        RECT  0.890 -0.300 1.110 0.340 ;
        RECT  1.110 -0.300 1.720 0.300 ;
        RECT  1.720 -0.300 1.940 0.340 ;
        RECT  1.940 -0.300 2.550 0.300 ;
        RECT  2.550 -0.300 2.770 0.340 ;
        RECT  2.770 -0.300 3.380 0.300 ;
        RECT  3.380 -0.300 3.600 0.340 ;
        RECT  3.600 -0.300 4.210 0.300 ;
        RECT  4.210 -0.300 4.430 0.340 ;
        RECT  4.430 -0.300 5.040 0.300 ;
        RECT  5.040 -0.300 5.260 0.340 ;
        RECT  5.260 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.620 2.820 ;
        RECT  0.620 2.180 0.840 2.820 ;
        RECT  0.840 2.220 1.420 2.820 ;
        RECT  1.420 2.180 1.640 2.820 ;
        RECT  1.640 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.580 1.630 2.800 2.050 ;
        RECT  2.040 1.930 2.580 2.050 ;
        RECT  1.820 1.370 2.040 2.050 ;
        RECT  1.240 1.930 1.820 2.050 ;
        RECT  3.720 1.370 3.940 1.790 ;
        RECT  3.180 1.370 3.720 1.490 ;
        RECT  2.960 1.370 3.180 2.050 ;
        RECT  2.420 1.370 2.960 1.490 ;
        RECT  4.860 1.630 5.080 2.050 ;
        RECT  4.320 1.930 4.860 2.050 ;
        RECT  4.100 1.370 4.320 2.050 ;
        RECT  3.560 1.930 4.100 2.050 ;
        RECT  3.340 1.630 3.560 2.050 ;
        RECT  2.200 1.370 2.420 1.790 ;
        RECT  1.020 1.370 1.240 2.050 ;
    END
END NR4D2

MACRO NR4D3
    CLASS CORE ;
    FOREIGN NR4D3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.600 1.370 6.670 1.790 ;
        RECT  0.150 0.470 6.670 0.630 ;
        RECT  6.670 0.470 6.820 1.790 ;
        RECT  6.820 0.470 7.090 1.490 ;
        RECT  7.090 1.370 7.360 1.490 ;
        RECT  7.360 1.370 7.580 1.790 ;
        RECT  7.580 1.370 8.120 1.490 ;
        RECT  8.120 1.370 8.340 2.050 ;
        RECT  7.090 0.470 8.710 0.630 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.830 1.530 1.235 ;
        RECT  1.530 1.005 1.830 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.830 3.450 1.235 ;
        RECT  3.450 1.005 3.750 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.830 5.370 1.235 ;
        RECT  5.370 1.005 5.670 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 0.830 7.610 1.235 ;
        RECT  7.610 1.005 7.910 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.590 0.300 ;
        RECT  0.590 -0.300 0.810 0.340 ;
        RECT  0.810 -0.300 1.420 0.300 ;
        RECT  1.420 -0.300 1.640 0.340 ;
        RECT  1.640 -0.300 2.250 0.300 ;
        RECT  2.250 -0.300 2.470 0.340 ;
        RECT  2.470 -0.300 3.080 0.300 ;
        RECT  3.080 -0.300 3.300 0.340 ;
        RECT  3.300 -0.300 3.910 0.300 ;
        RECT  3.910 -0.300 4.130 0.340 ;
        RECT  4.130 -0.300 4.740 0.300 ;
        RECT  4.740 -0.300 4.960 0.340 ;
        RECT  4.960 -0.300 5.570 0.300 ;
        RECT  5.570 -0.300 5.790 0.340 ;
        RECT  5.790 -0.300 6.400 0.300 ;
        RECT  6.400 -0.300 6.620 0.340 ;
        RECT  6.620 -0.300 7.220 0.300 ;
        RECT  7.220 -0.300 7.440 0.340 ;
        RECT  7.440 -0.300 8.050 0.300 ;
        RECT  8.050 -0.300 8.270 0.340 ;
        RECT  8.270 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.940 1.630 4.160 2.050 ;
        RECT  3.400 1.930 3.940 2.050 ;
        RECT  3.180 1.630 3.400 2.050 ;
        RECT  2.640 1.930 3.180 2.050 ;
        RECT  2.420 1.370 2.640 2.050 ;
        RECT  1.910 1.930 2.420 2.050 ;
        RECT  1.690 1.370 1.910 2.050 ;
        RECT  1.180 1.930 1.690 2.050 ;
        RECT  5.840 1.370 6.060 1.790 ;
        RECT  5.300 1.370 5.840 1.490 ;
        RECT  5.080 1.370 5.300 1.790 ;
        RECT  4.540 1.370 5.080 1.490 ;
        RECT  4.320 1.370 4.540 2.050 ;
        RECT  3.780 1.370 4.320 1.490 ;
        RECT  3.560 1.370 3.780 1.790 ;
        RECT  3.020 1.370 3.560 1.490 ;
        RECT  7.740 1.630 7.960 2.050 ;
        RECT  7.200 1.930 7.740 2.050 ;
        RECT  6.980 1.630 7.200 2.050 ;
        RECT  6.440 1.930 6.980 2.050 ;
        RECT  6.220 1.370 6.440 2.050 ;
        RECT  5.680 1.930 6.220 2.050 ;
        RECT  5.460 1.630 5.680 2.050 ;
        RECT  4.920 1.930 5.460 2.050 ;
        RECT  4.700 1.630 4.920 2.050 ;
        RECT  2.800 1.370 3.020 1.790 ;
        RECT  0.960 1.370 1.180 2.050 ;
        LAYER M1 ;
        RECT  8.120 1.370 8.340 2.050 ;
        RECT  7.580 1.370 8.120 1.490 ;
        RECT  7.360 1.370 7.580 1.790 ;
        RECT  0.150 0.470 6.455 0.630 ;
        RECT  7.305 0.470 8.710 0.630 ;
        RECT  7.305 1.370 7.360 1.490 ;
    END
END NR4D3

MACRO NR4D4
    CLASS CORE ;
    FOREIGN NR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.140 1.360 8.270 1.780 ;
        RECT  0.720 0.470 8.270 0.630 ;
        RECT  8.270 0.470 8.360 1.780 ;
        RECT  8.360 0.470 8.690 1.480 ;
        RECT  8.690 1.360 8.900 1.480 ;
        RECT  8.900 1.360 9.120 1.780 ;
        RECT  9.120 1.360 9.660 1.480 ;
        RECT  9.660 1.360 9.880 1.780 ;
        RECT  8.690 0.470 10.110 0.630 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.830 1.530 1.235 ;
        RECT  1.530 1.005 1.830 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 0.830 4.090 1.235 ;
        RECT  4.090 1.005 4.390 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.490 0.830 6.650 1.235 ;
        RECT  6.650 1.005 6.950 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.050 0.830 9.210 1.235 ;
        RECT  9.210 1.005 9.510 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.330 0.300 ;
        RECT  0.330 -0.300 0.550 0.340 ;
        RECT  0.550 -0.300 1.160 0.300 ;
        RECT  1.160 -0.300 1.380 0.340 ;
        RECT  1.380 -0.300 1.990 0.300 ;
        RECT  1.990 -0.300 2.210 0.340 ;
        RECT  2.210 -0.300 2.820 0.300 ;
        RECT  2.820 -0.300 3.040 0.340 ;
        RECT  3.040 -0.300 3.650 0.300 ;
        RECT  3.650 -0.300 3.870 0.340 ;
        RECT  3.870 -0.300 4.480 0.300 ;
        RECT  4.480 -0.300 4.700 0.340 ;
        RECT  4.700 -0.300 5.310 0.300 ;
        RECT  5.310 -0.300 5.530 0.340 ;
        RECT  5.530 -0.300 6.140 0.300 ;
        RECT  6.140 -0.300 6.360 0.340 ;
        RECT  6.360 -0.300 6.970 0.300 ;
        RECT  6.970 -0.300 7.190 0.340 ;
        RECT  7.190 -0.300 7.800 0.300 ;
        RECT  7.800 -0.300 8.020 0.340 ;
        RECT  8.020 -0.300 8.620 0.300 ;
        RECT  8.620 -0.300 8.840 0.340 ;
        RECT  8.840 -0.300 9.450 0.300 ;
        RECT  9.450 -0.300 9.670 0.340 ;
        RECT  9.670 -0.300 10.280 0.300 ;
        RECT  10.280 -0.300 10.500 0.340 ;
        RECT  10.500 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.120 1.620 5.340 2.040 ;
        RECT  4.580 1.920 5.120 2.040 ;
        RECT  4.360 1.620 4.580 2.040 ;
        RECT  3.820 1.920 4.360 2.040 ;
        RECT  3.600 1.620 3.820 2.040 ;
        RECT  3.060 1.920 3.600 2.040 ;
        RECT  2.840 1.360 3.060 2.040 ;
        RECT  2.320 1.920 2.840 2.040 ;
        RECT  2.100 1.360 2.320 2.040 ;
        RECT  1.580 1.920 2.100 2.040 ;
        RECT  1.360 1.360 1.580 2.040 ;
        RECT  0.840 1.920 1.360 2.040 ;
        RECT  7.380 1.360 7.600 1.780 ;
        RECT  6.840 1.360 7.380 1.480 ;
        RECT  6.620 1.360 6.840 1.780 ;
        RECT  6.080 1.360 6.620 1.480 ;
        RECT  5.860 1.360 6.080 1.780 ;
        RECT  4.960 1.360 5.860 1.480 ;
        RECT  4.740 1.360 4.960 1.780 ;
        RECT  4.200 1.360 4.740 1.480 ;
        RECT  3.980 1.360 4.200 1.780 ;
        RECT  3.440 1.360 3.980 1.480 ;
        RECT  10.040 1.360 10.260 2.040 ;
        RECT  9.500 1.900 10.040 2.040 ;
        RECT  9.280 1.620 9.500 2.040 ;
        RECT  8.740 1.900 9.280 2.040 ;
        RECT  8.520 1.620 8.740 2.040 ;
        RECT  7.980 1.900 8.520 2.040 ;
        RECT  7.760 1.620 7.980 2.040 ;
        RECT  7.220 1.900 7.760 2.040 ;
        RECT  7.000 1.620 7.220 2.040 ;
        RECT  6.460 1.900 7.000 2.040 ;
        RECT  6.240 1.620 6.460 2.040 ;
        RECT  5.700 1.900 6.240 2.040 ;
        RECT  5.480 1.620 5.700 2.040 ;
        RECT  3.220 1.360 3.440 1.780 ;
        RECT  0.620 1.360 0.840 2.040 ;
        LAYER M1 ;
        RECT  9.660 1.360 9.880 1.780 ;
        RECT  9.120 1.360 9.660 1.480 ;
        RECT  0.720 0.470 8.055 0.630 ;
        RECT  8.905 0.470 10.110 0.630 ;
        RECT  8.905 1.360 9.120 1.780 ;
    END
END NR4D4

MACRO NR4D8
    CLASS CORE ;
    FOREIGN NR4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.640 2.510 2.020 ;
        RECT  1.780 0.710 2.510 0.870 ;
        RECT  2.510 0.710 2.930 2.020 ;
        RECT  2.930 1.640 4.120 2.020 ;
        RECT  2.930 0.710 4.140 0.870 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 0.810 0.730 1.125 ;
        RECT  0.730 0.810 0.830 1.515 ;
        RECT  0.830 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.230 1.235 ;
        RECT  0.230 1.010 0.300 1.235 ;
        END
    END A1
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A4
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.295 0.300 ;
        RECT  4.295 -0.300 4.515 0.340 ;
        RECT  4.515 -0.300 5.085 0.300 ;
        RECT  5.085 -0.300 5.305 0.340 ;
        RECT  5.305 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 4.295 2.820 ;
        RECT  4.295 2.180 4.515 2.820 ;
        RECT  4.515 2.220 5.085 2.820 ;
        RECT  5.085 2.180 5.305 2.820 ;
        RECT  5.305 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.570 1.080 4.760 1.240 ;
        RECT  4.450 0.470 4.570 1.240 ;
        RECT  1.330 0.470 4.450 0.590 ;
        RECT  0.540 0.470 1.330 0.630 ;
        RECT  0.430 0.470 0.540 1.510 ;
        RECT  0.430 1.960 0.460 2.100 ;
        RECT  0.420 0.470 0.430 2.100 ;
        RECT  0.270 1.390 0.420 2.100 ;
        RECT  5.480 0.430 5.700 0.850 ;
        RECT  5.670 1.960 5.700 2.100 ;
        RECT  5.510 1.390 5.670 2.100 ;
        RECT  5.000 1.390 5.510 1.510 ;
        RECT  5.480 1.960 5.510 2.100 ;
        RECT  5.000 0.690 5.480 0.850 ;
        RECT  4.910 0.690 5.000 1.510 ;
        RECT  4.880 0.430 4.910 1.510 ;
        RECT  4.880 1.960 4.910 2.100 ;
        RECT  4.690 0.430 4.880 0.850 ;
        RECT  4.720 1.390 4.880 2.100 ;
        RECT  4.210 1.390 4.720 1.510 ;
        RECT  4.690 1.960 4.720 2.100 ;
        RECT  4.090 1.080 4.210 1.510 ;
        RECT  0.240 1.960 0.270 2.100 ;
        RECT  3.370 1.080 4.090 1.240 ;
        LAYER M1 ;
        RECT  1.780 0.710 2.295 0.870 ;
        RECT  1.800 1.640 2.295 2.020 ;
        RECT  3.145 0.710 4.140 0.870 ;
        RECT  3.145 1.640 4.120 2.020 ;
    END
END NR4D8

MACRO OA211D0
    CLASS CORE ;
    FOREIGN OA211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.660 2.150 2.090 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.080 0.790 1.240 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.910 1.080 1.050 1.240 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.670 0.300 ;
        RECT  1.670 -0.300 1.890 0.340 ;
        RECT  1.890 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.480 2.820 ;
        RECT  0.480 2.180 0.700 2.820 ;
        RECT  0.700 2.220 1.550 2.820 ;
        RECT  1.550 2.180 1.770 2.820 ;
        RECT  1.770 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.710 0.710 1.870 2.050 ;
        RECT  1.000 0.710 1.710 0.870 ;
        RECT  0.070 1.890 1.710 2.050 ;
    END
END OA211D0

MACRO OA211D1
    CLASS CORE ;
    FOREIGN OA211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.960 2.310 2.100 ;
        RECT  2.310 0.420 2.470 2.100 ;
        RECT  2.470 1.960 2.500 2.100 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 1.890 0.300 ;
        RECT  1.890 -0.300 2.110 0.340 ;
        RECT  2.110 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.490 2.820 ;
        RECT  1.490 2.180 1.710 2.820 ;
        RECT  1.710 2.220 1.890 2.820 ;
        RECT  1.890 2.180 2.110 2.820 ;
        RECT  2.110 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.450 1.770 0.610 ;
        RECT  0.990 0.470 1.530 0.610 ;
        RECT  2.030 0.730 2.190 1.770 ;
        RECT  1.130 0.730 2.030 0.885 ;
        RECT  1.070 1.650 2.030 1.770 ;
        RECT  0.850 1.650 1.070 2.070 ;
        RECT  0.250 1.650 0.850 1.770 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.090 1.370 0.250 2.100 ;
        RECT  0.770 0.470 0.990 0.885 ;
        RECT  0.060 1.960 0.090 2.100 ;
    END
END OA211D1

MACRO OA211D2
    CLASS CORE ;
    FOREIGN OA211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.960 2.270 2.100 ;
        RECT  2.270 1.390 2.330 2.100 ;
        RECT  2.270 0.420 2.330 0.900 ;
        RECT  2.330 0.420 2.430 2.100 ;
        RECT  2.430 1.960 2.460 2.100 ;
        RECT  2.430 0.780 2.470 1.515 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.180 0.680 2.820 ;
        RECT  0.680 2.220 1.490 2.820 ;
        RECT  1.490 2.180 1.710 2.820 ;
        RECT  1.710 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.530 0.450 1.770 0.610 ;
        RECT  0.990 0.470 1.530 0.610 ;
        RECT  2.110 1.080 2.210 1.240 ;
        RECT  1.990 0.730 2.110 1.770 ;
        RECT  1.130 0.730 1.990 0.885 ;
        RECT  1.070 1.650 1.990 1.770 ;
        RECT  0.850 1.650 1.070 2.070 ;
        RECT  0.250 1.650 0.850 1.770 ;
        RECT  0.250 1.960 0.280 2.100 ;
        RECT  0.090 1.370 0.250 2.100 ;
        RECT  0.060 1.960 0.090 2.100 ;
        RECT  0.770 0.470 0.990 0.885 ;
    END
END OA211D2

MACRO OA211D4
    CLASS CORE ;
    FOREIGN OA211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.650 3.790 2.030 ;
        RECT  3.610 0.490 3.790 0.870 ;
        RECT  3.790 0.490 4.210 2.030 ;
        RECT  4.210 1.650 4.610 2.030 ;
        RECT  4.210 0.490 4.610 0.870 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.755 ;
        RECT  0.250 1.635 1.230 1.755 ;
        RECT  1.230 1.030 1.390 1.755 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.660 1.030 1.820 1.755 ;
        RECT  1.820 1.635 2.650 1.755 ;
        RECT  2.650 1.005 2.770 1.755 ;
        RECT  2.770 1.005 3.110 1.235 ;
        END
    END A1
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END C
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.700 0.300 ;
        RECT  0.700 -0.300 0.920 0.340 ;
        RECT  0.920 -0.300 3.220 0.300 ;
        RECT  3.220 -0.300 3.440 0.340 ;
        RECT  3.440 -0.300 4.000 0.300 ;
        RECT  4.000 -0.300 4.220 0.340 ;
        RECT  4.220 -0.300 4.780 0.300 ;
        RECT  4.780 -0.300 5.000 0.340 ;
        RECT  5.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.770 2.820 ;
        RECT  2.770 2.190 2.990 2.820 ;
        RECT  2.990 2.220 3.210 2.820 ;
        RECT  3.210 2.180 3.430 2.820 ;
        RECT  3.430 2.220 4.000 2.820 ;
        RECT  4.000 2.190 4.220 2.820 ;
        RECT  4.220 2.220 4.780 2.820 ;
        RECT  4.780 2.190 5.000 2.820 ;
        RECT  5.000 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.870 0.440 3.110 0.600 ;
        RECT  2.330 0.470 2.870 0.600 ;
        RECT  2.110 0.440 2.330 0.600 ;
        RECT  1.570 0.470 2.110 0.600 ;
        RECT  1.350 0.470 1.570 0.890 ;
        RECT  0.280 0.470 1.350 0.630 ;
        RECT  3.240 0.720 3.400 2.050 ;
        RECT  1.710 0.720 3.240 0.880 ;
        RECT  0.400 1.890 3.240 2.050 ;
        RECT  0.060 0.470 0.280 0.885 ;
        LAYER M1 ;
        RECT  4.425 0.490 4.610 0.870 ;
        RECT  4.425 1.650 4.610 2.030 ;
    END
END OA211D4

MACRO OA21D0
    CLASS CORE ;
    FOREIGN OA21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.660 1.830 2.090 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.240 0.300 ;
        RECT  1.240 -0.300 1.460 0.340 ;
        RECT  1.460 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.230 2.820 ;
        RECT  1.230 2.180 1.450 2.820 ;
        RECT  1.450 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.470 1.020 0.880 ;
        RECT  0.260 0.470 0.860 0.590 ;
        RECT  1.390 1.030 1.550 2.050 ;
        RECT  0.570 1.890 1.390 2.050 ;
        RECT  0.450 0.710 0.570 2.050 ;
        RECT  0.100 0.470 0.260 0.880 ;
        RECT  0.570 0.710 0.690 0.870 ;
    END
END OA21D0

MACRO OA21D1
    CLASS CORE ;
    FOREIGN OA21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.670 0.420 1.830 2.100 ;
        RECT  1.830 1.960 1.860 2.100 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.240 0.300 ;
        RECT  1.240 -0.300 1.460 0.340 ;
        RECT  1.460 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.230 2.820 ;
        RECT  1.230 2.180 1.450 2.820 ;
        RECT  1.450 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.470 1.020 0.880 ;
        RECT  0.260 0.470 0.860 0.590 ;
        RECT  1.360 1.030 1.520 1.760 ;
        RECT  1.030 1.640 1.360 1.760 ;
        RECT  0.810 1.640 1.030 2.060 ;
        RECT  0.570 1.640 0.810 1.760 ;
        RECT  0.570 0.710 0.690 0.870 ;
        RECT  0.100 0.470 0.260 0.880 ;
        RECT  0.450 0.710 0.570 1.760 ;
    END
END OA21D1

MACRO OA21D2
    CLASS CORE ;
    FOREIGN OA21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.960 1.630 2.100 ;
        RECT  1.630 1.390 1.690 2.100 ;
        RECT  1.630 0.420 1.690 0.900 ;
        RECT  1.690 0.420 1.790 2.100 ;
        RECT  1.790 1.960 1.820 2.100 ;
        RECT  1.790 0.780 1.830 1.515 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.210 2.820 ;
        RECT  1.210 2.180 1.430 2.820 ;
        RECT  1.430 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.860 0.470 1.020 0.880 ;
        RECT  0.260 0.470 0.860 0.590 ;
        RECT  1.350 1.030 1.510 1.760 ;
        RECT  1.030 1.640 1.350 1.760 ;
        RECT  0.810 1.640 1.030 2.060 ;
        RECT  0.570 1.640 0.810 1.760 ;
        RECT  0.570 0.710 0.690 0.870 ;
        RECT  0.450 0.710 0.570 1.760 ;
        RECT  0.100 0.470 0.260 0.880 ;
    END
END OA21D2

MACRO OA21D4
    CLASS CORE ;
    FOREIGN OA21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.650 3.150 2.030 ;
        RECT  2.630 0.490 3.150 0.870 ;
        RECT  3.150 0.490 3.570 2.030 ;
        RECT  3.570 1.650 3.640 2.030 ;
        RECT  3.570 0.490 3.640 0.870 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.250 1.080 0.410 1.240 ;
        RECT  0.410 1.005 0.550 1.755 ;
        RECT  0.550 1.635 2.100 1.755 ;
        RECT  2.100 1.030 2.260 1.755 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.030 0.840 1.515 ;
        RECT  0.840 1.395 1.690 1.515 ;
        RECT  1.690 1.035 1.830 1.515 ;
        RECT  1.830 1.080 1.950 1.240 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.020 0.300 ;
        RECT  3.020 -0.300 3.240 0.340 ;
        RECT  3.240 -0.300 3.810 0.300 ;
        RECT  3.810 -0.300 4.030 0.340 ;
        RECT  4.030 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.180 2.820 ;
        RECT  1.180 2.180 1.400 2.820 ;
        RECT  1.400 2.220 2.240 2.820 ;
        RECT  2.240 2.180 2.460 2.820 ;
        RECT  2.460 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 3.810 2.820 ;
        RECT  3.810 2.180 4.030 2.820 ;
        RECT  4.030 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.940 0.440 2.180 0.600 ;
        RECT  1.400 0.470 1.940 0.600 ;
        RECT  1.180 0.440 1.400 0.600 ;
        RECT  0.640 0.470 1.180 0.600 ;
        RECT  2.510 1.080 2.740 1.240 ;
        RECT  2.390 0.720 2.510 2.050 ;
        RECT  0.780 0.720 2.390 0.880 ;
        RECT  0.420 0.470 0.640 0.885 ;
        RECT  0.500 1.890 2.390 2.050 ;
        LAYER M1 ;
        RECT  2.630 0.490 2.935 0.870 ;
        RECT  2.630 1.650 2.935 2.030 ;
    END
END OA21D4

MACRO OA221D0
    CLASS CORE ;
    FOREIGN OA221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.570 2.470 2.070 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.285 1.850 1.795 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.140 1.530 1.795 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.755 ;
        RECT  0.250 1.635 1.090 1.755 ;
        RECT  1.090 1.480 1.250 1.755 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.190 1.050 1.350 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.870 0.300 ;
        RECT  1.870 -0.300 2.090 0.350 ;
        RECT  2.090 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.910 2.820 ;
        RECT  0.910 2.180 1.130 2.820 ;
        RECT  1.130 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.070 0.660 0.500 0.820 ;
        RECT  0.220 1.890 0.460 2.050 ;
        RECT  0.740 0.710 1.210 0.870 ;
        RECT  1.210 0.710 1.330 1.020 ;
        RECT  0.460 1.915 2.020 2.050 ;
        RECT  1.330 0.900 2.020 1.020 ;
        RECT  2.020 0.900 2.180 2.050 ;
        RECT  0.500 0.470 0.620 0.820 ;
        RECT  0.620 0.470 1.450 0.590 ;
        RECT  1.450 0.470 1.670 0.780 ;
    END
END OA221D0

MACRO OA221D1
    CLASS CORE ;
    FOREIGN OA221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.060 2.170 1.795 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.190 2.820 ;
        RECT  0.190 2.180 0.410 2.820 ;
        RECT  0.410 2.220 1.500 2.820 ;
        RECT  1.500 2.180 1.720 2.820 ;
        RECT  1.720 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 1.030 2.470 2.050 ;
        RECT  2.470 1.030 2.510 1.270 ;
        RECT  1.890 0.720 2.050 0.940 ;
        RECT  0.300 0.470 0.840 0.590 ;
        RECT  0.840 0.470 1.060 0.885 ;
        RECT  1.060 0.470 1.600 0.590 ;
        RECT  1.600 0.420 1.840 0.590 ;
        RECT  2.080 1.930 2.350 2.050 ;
        RECT  1.860 1.930 2.080 2.090 ;
        RECT  1.070 1.930 1.860 2.050 ;
        RECT  0.850 1.635 1.070 2.050 ;
        RECT  0.280 1.635 0.850 1.755 ;
        RECT  0.280 0.710 0.700 0.870 ;
        RECT  1.200 0.720 1.890 0.880 ;
        RECT  0.060 0.430 0.300 0.590 ;
        RECT  0.160 0.710 0.280 1.755 ;
    END
END OA221D1

MACRO OA221D2
    CLASS CORE ;
    FOREIGN OA221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.960 2.590 2.100 ;
        RECT  2.590 1.390 2.650 2.100 ;
        RECT  2.590 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.750 2.100 ;
        RECT  2.750 1.960 2.780 2.100 ;
        RECT  2.750 0.780 2.790 1.515 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.060 2.170 1.795 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.190 2.820 ;
        RECT  0.190 2.180 0.410 2.820 ;
        RECT  0.410 2.220 1.500 2.820 ;
        RECT  1.500 2.180 1.720 2.820 ;
        RECT  1.720 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.600 0.420 1.840 0.590 ;
        RECT  1.060 0.470 1.600 0.590 ;
        RECT  0.840 0.470 1.060 0.885 ;
        RECT  0.300 0.470 0.840 0.590 ;
        RECT  1.890 0.720 2.050 0.940 ;
        RECT  2.440 1.050 2.520 1.270 ;
        RECT  2.320 1.050 2.440 2.050 ;
        RECT  2.080 1.930 2.320 2.050 ;
        RECT  1.860 1.930 2.080 2.090 ;
        RECT  1.070 1.930 1.860 2.050 ;
        RECT  0.850 1.635 1.070 2.050 ;
        RECT  0.280 1.635 0.850 1.755 ;
        RECT  0.280 0.710 0.700 0.870 ;
        RECT  0.160 0.710 0.280 1.755 ;
        RECT  1.200 0.720 1.890 0.880 ;
        RECT  0.060 0.430 0.300 0.590 ;
    END
END OA221D2

MACRO OA221D4
    CLASS CORE ;
    FOREIGN OA221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.800 1.650 5.070 2.030 ;
        RECT  4.800 0.490 5.070 0.870 ;
        RECT  5.070 0.490 5.490 2.030 ;
        RECT  5.490 1.650 5.840 2.030 ;
        RECT  5.490 0.490 5.840 0.870 ;
        END
    END Z
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.030 1.220 1.475 ;
        RECT  1.220 1.355 2.010 1.475 ;
        RECT  2.010 1.005 2.130 1.475 ;
        RECT  2.130 1.005 2.470 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 2.990 1.235 ;
        RECT  2.990 1.005 3.110 1.475 ;
        RECT  3.110 1.355 3.920 1.475 ;
        RECT  3.920 1.030 4.080 1.475 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.210 0.300 ;
        RECT  5.210 -0.300 5.430 0.340 ;
        RECT  5.430 -0.300 6.030 0.300 ;
        RECT  6.030 -0.300 6.250 0.340 ;
        RECT  6.250 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.490 2.820 ;
        RECT  0.490 2.180 0.710 2.820 ;
        RECT  0.710 2.220 1.570 2.820 ;
        RECT  1.570 2.180 1.790 2.820 ;
        RECT  1.790 2.220 3.360 2.820 ;
        RECT  3.360 2.180 3.580 2.820 ;
        RECT  3.580 2.220 4.390 2.820 ;
        RECT  4.390 2.180 4.610 2.820 ;
        RECT  4.610 2.220 5.210 2.820 ;
        RECT  5.210 2.180 5.430 2.820 ;
        RECT  5.430 2.220 6.030 2.820 ;
        RECT  6.030 2.180 6.250 2.820 ;
        RECT  6.250 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.990 0.470 2.510 0.620 ;
        RECT  0.770 0.470 0.990 0.890 ;
        RECT  0.290 0.470 0.770 0.610 ;
        RECT  4.520 0.770 4.680 1.750 ;
        RECT  4.370 0.770 4.520 0.890 ;
        RECT  4.240 1.630 4.520 1.750 ;
        RECT  4.150 0.470 4.370 0.890 ;
        RECT  4.020 1.630 4.240 2.050 ;
        RECT  2.630 0.470 4.150 0.620 ;
        RECT  2.910 1.910 4.020 2.050 ;
        RECT  2.870 1.910 2.910 2.100 ;
        RECT  2.720 1.370 2.870 2.100 ;
        RECT  2.690 1.910 2.720 2.100 ;
        RECT  2.450 1.910 2.690 2.050 ;
        RECT  2.420 1.910 2.450 2.100 ;
        RECT  2.260 1.370 2.420 2.100 ;
        RECT  2.230 1.910 2.260 2.100 ;
        RECT  1.120 1.910 2.230 2.050 ;
        RECT  0.900 1.630 1.120 2.050 ;
        RECT  0.290 1.910 0.900 2.050 ;
        RECT  0.260 1.910 0.290 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  1.130 0.740 4.010 0.885 ;
        RECT  0.070 0.470 0.290 0.890 ;
        RECT  0.070 1.960 0.100 2.100 ;
        LAYER M1 ;
        RECT  4.800 0.490 4.855 0.870 ;
        RECT  4.800 1.650 4.855 2.030 ;
        RECT  5.700 0.490 5.840 0.870 ;
        RECT  5.705 1.650 5.840 2.030 ;
    END
END OA221D4

MACRO OA222D0
    CLASS CORE ;
    FOREIGN OA222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 0.660 3.110 1.710 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.080 0.390 1.240 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.490 1.490 1.760 ;
        RECT  1.490 1.640 2.310 1.760 ;
        RECT  2.310 1.005 2.470 1.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.540 1.200 1.690 1.360 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.430 0.300 ;
        RECT  0.430 -0.300 0.650 0.340 ;
        RECT  0.650 -0.300 2.630 0.300 ;
        RECT  2.630 -0.300 2.850 0.340 ;
        RECT  2.850 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.470 2.820 ;
        RECT  1.470 2.180 1.690 2.820 ;
        RECT  1.690 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.280 0.430 2.520 0.590 ;
        RECT  1.140 0.470 2.280 0.590 ;
        RECT  1.020 0.470 1.140 0.820 ;
        RECT  2.670 0.710 2.830 2.050 ;
        RECT  1.510 0.710 2.670 0.870 ;
        RECT  0.780 1.890 2.670 2.050 ;
        RECT  0.070 0.660 1.020 0.820 ;
    END
END OA222D0

MACRO OA222D1
    CLASS CORE ;
    FOREIGN OA222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.960 2.950 2.100 ;
        RECT  2.950 1.390 2.980 2.100 ;
        RECT  2.950 0.420 2.980 0.955 ;
        RECT  2.980 0.420 3.110 2.100 ;
        RECT  3.110 1.960 3.140 2.100 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.580 1.240 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.170 2.820 ;
        RECT  0.170 2.180 0.390 2.820 ;
        RECT  0.390 2.220 1.500 2.820 ;
        RECT  1.500 2.180 1.720 2.820 ;
        RECT  1.720 2.220 2.520 2.820 ;
        RECT  2.520 2.180 2.740 2.820 ;
        RECT  2.740 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.860 1.640 2.080 2.060 ;
        RECT  2.080 1.640 2.700 1.760 ;
        RECT  2.700 1.050 2.820 1.760 ;
        RECT  2.820 1.050 2.860 1.270 ;
        RECT  2.220 0.450 2.440 0.870 ;
        RECT  0.280 0.470 0.820 0.590 ;
        RECT  0.820 0.470 1.040 0.885 ;
        RECT  1.040 0.470 1.580 0.590 ;
        RECT  1.580 0.430 1.820 0.590 ;
        RECT  1.060 1.640 1.860 1.760 ;
        RECT  0.840 1.640 1.060 2.060 ;
        RECT  0.260 1.640 0.840 1.760 ;
        RECT  0.260 0.710 0.680 0.870 ;
        RECT  1.180 0.710 2.220 0.870 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.140 0.710 0.260 1.760 ;
    END
END OA222D1

MACRO OA222D2
    CLASS CORE ;
    FOREIGN OA222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.960 2.950 2.100 ;
        RECT  2.950 1.390 2.980 2.100 ;
        RECT  2.950 0.420 2.980 0.955 ;
        RECT  2.980 0.420 3.110 2.100 ;
        RECT  3.110 1.960 3.140 2.100 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.080 2.580 1.240 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.335 0.300 ;
        RECT  3.335 -0.300 3.555 0.340 ;
        RECT  3.555 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.170 2.820 ;
        RECT  0.170 2.180 0.390 2.820 ;
        RECT  0.390 2.220 1.500 2.820 ;
        RECT  1.500 2.180 1.720 2.820 ;
        RECT  1.720 2.220 2.520 2.820 ;
        RECT  2.520 2.180 2.740 2.820 ;
        RECT  2.740 2.220 3.335 2.820 ;
        RECT  3.335 2.180 3.555 2.820 ;
        RECT  3.555 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.580 0.430 1.820 0.590 ;
        RECT  1.040 0.470 1.580 0.590 ;
        RECT  0.820 0.470 1.040 0.885 ;
        RECT  0.280 0.470 0.820 0.590 ;
        RECT  2.220 0.450 2.440 0.870 ;
        RECT  2.820 1.050 2.860 1.270 ;
        RECT  2.700 1.050 2.820 1.760 ;
        RECT  2.080 1.640 2.700 1.760 ;
        RECT  1.860 1.640 2.080 2.060 ;
        RECT  1.060 1.640 1.860 1.760 ;
        RECT  0.840 1.640 1.060 2.060 ;
        RECT  0.260 1.640 0.840 1.760 ;
        RECT  0.260 0.710 0.680 0.870 ;
        RECT  0.140 0.710 0.260 1.760 ;
        RECT  1.180 0.710 2.220 0.870 ;
        RECT  0.060 0.430 0.280 0.590 ;
    END
END OA222D2

MACRO OA222D4
    CLASS CORE ;
    FOREIGN OA222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.630 1.650 6.030 2.030 ;
        RECT  5.630 0.490 6.030 0.870 ;
        RECT  6.030 0.490 6.450 2.030 ;
        RECT  6.450 1.650 6.580 2.030 ;
        RECT  6.450 0.490 6.580 0.870 ;
        END
    END Z
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.395 1.380 1.515 ;
        RECT  1.380 1.030 1.540 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.515 ;
        RECT  2.150 1.395 2.910 1.515 ;
        RECT  2.910 1.030 3.070 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.630 1.235 ;
        RECT  3.630 1.005 3.750 1.515 ;
        RECT  3.750 1.395 4.700 1.515 ;
        RECT  4.700 1.030 4.860 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.210 2.820 ;
        RECT  0.210 2.180 0.430 2.820 ;
        RECT  0.430 2.220 1.530 2.820 ;
        RECT  1.530 2.180 1.750 2.820 ;
        RECT  1.750 2.220 2.980 2.820 ;
        RECT  2.980 2.180 3.200 2.820 ;
        RECT  3.200 2.220 4.150 2.820 ;
        RECT  4.150 2.180 4.370 2.820 ;
        RECT  4.370 2.220 5.220 2.820 ;
        RECT  5.220 2.180 5.440 2.820 ;
        RECT  5.440 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.790 0.725 3.310 0.885 ;
        RECT  1.570 0.465 1.790 0.885 ;
        RECT  1.090 0.725 1.570 0.885 ;
        RECT  0.870 0.465 1.090 0.885 ;
        RECT  0.290 0.725 0.870 0.885 ;
        RECT  4.570 0.445 4.810 0.605 ;
        RECT  4.030 0.485 4.570 0.605 ;
        RECT  3.810 0.445 4.030 0.605 ;
        RECT  2.930 0.485 3.810 0.605 ;
        RECT  2.710 0.445 2.930 0.605 ;
        RECT  2.170 0.485 2.710 0.605 ;
        RECT  5.315 0.725 5.475 1.755 ;
        RECT  5.170 0.725 5.315 0.885 ;
        RECT  5.040 1.635 5.315 1.755 ;
        RECT  4.950 0.465 5.170 0.885 ;
        RECT  4.820 1.635 5.040 2.050 ;
        RECT  3.430 0.725 4.950 0.885 ;
        RECT  3.710 1.635 4.820 1.755 ;
        RECT  3.490 1.635 3.710 2.050 ;
        RECT  2.420 1.635 3.490 1.755 ;
        RECT  2.200 1.635 2.420 2.050 ;
        RECT  1.090 1.635 2.200 1.755 ;
        RECT  0.870 1.635 1.090 2.050 ;
        RECT  1.930 0.445 2.170 0.605 ;
        RECT  0.070 0.465 0.290 0.885 ;
        LAYER M1 ;
        RECT  5.630 0.490 5.815 0.870 ;
        RECT  5.630 1.650 5.815 2.030 ;
    END
END OA222D4

MACRO OA22D0
    CLASS CORE ;
    FOREIGN OA22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.430 2.150 2.030 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.370 0.700 1.795 ;
        RECT  0.700 1.675 1.370 1.795 ;
        RECT  1.370 1.005 1.510 1.795 ;
        RECT  1.510 1.360 1.600 1.580 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.110 1.250 1.330 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.985 0.250 1.515 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.460 2.820 ;
        RECT  1.460 2.180 1.680 2.820 ;
        RECT  1.680 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.660 0.470 1.220 0.590 ;
        RECT  1.220 0.430 1.460 0.590 ;
        RECT  1.720 0.710 1.870 2.035 ;
        RECT  0.810 0.710 1.720 0.870 ;
        RECT  0.930 1.915 1.720 2.035 ;
        RECT  0.690 1.915 0.930 2.075 ;
        RECT  0.420 0.430 0.660 0.590 ;
    END
END OA22D0

MACRO OA22D1
    CLASS CORE ;
    FOREIGN OA22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.960 2.310 2.100 ;
        RECT  2.310 0.420 2.470 2.100 ;
        RECT  2.470 1.960 2.500 2.100 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.890 0.300 ;
        RECT  1.890 -0.300 2.110 0.340 ;
        RECT  2.110 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.800 2.820 ;
        RECT  0.800 2.180 1.020 2.820 ;
        RECT  1.020 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.450 1.780 0.610 ;
        RECT  1.000 0.470 1.540 0.610 ;
        RECT  0.780 0.470 1.000 0.885 ;
        RECT  0.280 0.470 0.780 0.610 ;
        RECT  1.980 0.730 2.140 1.760 ;
        RECT  1.140 0.730 1.980 0.885 ;
        RECT  1.690 1.640 1.980 1.760 ;
        RECT  1.470 1.640 1.690 2.060 ;
        RECT  0.360 1.640 1.470 1.760 ;
        RECT  0.140 1.640 0.360 2.060 ;
        RECT  0.060 0.470 0.280 0.885 ;
    END
END OA22D1

MACRO OA22D2
    CLASS CORE ;
    FOREIGN OA22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.240 1.960 2.270 2.100 ;
        RECT  2.270 1.390 2.330 2.100 ;
        RECT  2.270 0.420 2.330 0.900 ;
        RECT  2.330 0.420 2.430 2.100 ;
        RECT  2.430 1.960 2.460 2.100 ;
        RECT  2.430 0.780 2.470 1.515 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.800 2.820 ;
        RECT  0.800 2.180 1.020 2.820 ;
        RECT  1.020 2.220 1.850 2.820 ;
        RECT  1.850 2.180 2.070 2.820 ;
        RECT  2.070 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.450 1.780 0.610 ;
        RECT  1.000 0.470 1.540 0.610 ;
        RECT  0.780 0.470 1.000 0.885 ;
        RECT  0.280 0.470 0.780 0.610 ;
        RECT  1.990 0.730 2.150 1.760 ;
        RECT  1.140 0.730 1.990 0.885 ;
        RECT  1.690 1.640 1.990 1.760 ;
        RECT  1.470 1.640 1.690 2.060 ;
        RECT  0.360 1.640 1.470 1.760 ;
        RECT  0.060 0.470 0.280 0.885 ;
        RECT  0.140 1.640 0.360 2.060 ;
    END
END OA22D2

MACRO OA22D4
    CLASS CORE ;
    FOREIGN OA22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.650 4.110 2.030 ;
        RECT  3.750 0.490 4.110 0.870 ;
        RECT  4.110 0.490 4.530 2.030 ;
        RECT  4.530 1.650 4.680 2.030 ;
        RECT  4.530 0.490 4.680 0.870 ;
        END
    END Z
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.475 ;
        RECT  2.150 1.355 2.910 1.475 ;
        RECT  2.910 1.030 3.070 1.475 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        RECT  0.570 1.395 1.390 1.515 ;
        RECT  1.390 1.030 1.550 1.515 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.340 ;
        RECT  0.690 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.220 2.820 ;
        RECT  0.220 2.180 0.440 2.820 ;
        RECT  0.440 2.220 1.600 2.820 ;
        RECT  1.600 2.180 1.820 2.820 ;
        RECT  1.820 2.220 2.970 2.820 ;
        RECT  2.970 2.180 3.190 2.820 ;
        RECT  3.190 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.090 0.440 3.330 0.600 ;
        RECT  2.550 0.470 3.090 0.600 ;
        RECT  2.330 0.440 2.550 0.600 ;
        RECT  1.790 0.470 2.330 0.600 ;
        RECT  1.570 0.470 1.790 0.885 ;
        RECT  1.100 0.470 1.570 0.590 ;
        RECT  0.880 0.470 1.100 0.885 ;
        RECT  0.280 0.470 0.880 0.590 ;
        RECT  3.435 0.720 3.595 1.755 ;
        RECT  1.930 0.720 3.435 0.880 ;
        RECT  2.550 1.635 3.435 1.755 ;
        RECT  2.330 1.635 2.550 2.050 ;
        RECT  1.100 1.635 2.330 1.755 ;
        RECT  0.060 0.470 0.280 0.890 ;
        RECT  0.880 1.635 1.100 2.050 ;
        LAYER M1 ;
        RECT  3.750 0.490 3.895 0.870 ;
        RECT  3.750 1.650 3.895 2.030 ;
    END
END OA22D4

MACRO OA31D0
    CLASS CORE ;
    FOREIGN OA31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.660 2.150 1.990 ;
        END
    END Z
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 1.490 2.820 ;
        RECT  1.490 2.180 1.710 2.820 ;
        RECT  1.710 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.715 0.710 1.870 1.940 ;
        RECT  0.070 0.710 1.715 0.870 ;
        RECT  1.050 1.780 1.715 1.940 ;
    END
END OA31D0

MACRO OA31D1
    CLASS CORE ;
    FOREIGN OA31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  1.990 0.420 2.150 2.100 ;
        RECT  2.150 1.960 2.180 2.100 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.540 2.820 ;
        RECT  1.540 2.180 1.760 2.820 ;
        RECT  1.760 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.440 1.450 0.600 ;
        RECT  0.670 0.470 1.210 0.600 ;
        RECT  1.710 0.720 1.870 1.755 ;
        RECT  0.290 0.720 1.710 0.880 ;
        RECT  1.340 1.635 1.710 1.755 ;
        RECT  1.120 1.635 1.340 2.050 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.430 0.440 0.670 0.600 ;
    END
END OA31D1

MACRO OA31D2
    CLASS CORE ;
    FOREIGN OA31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.950 1.390 2.010 2.100 ;
        RECT  1.950 0.420 2.010 0.900 ;
        RECT  2.010 0.420 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.780 2.150 1.515 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.520 2.820 ;
        RECT  1.520 2.180 1.740 2.820 ;
        RECT  1.740 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.440 1.450 0.600 ;
        RECT  0.670 0.470 1.210 0.600 ;
        RECT  1.830 1.050 1.880 1.270 ;
        RECT  1.710 0.720 1.830 1.755 ;
        RECT  0.290 0.720 1.710 0.880 ;
        RECT  1.340 1.635 1.710 1.755 ;
        RECT  1.120 1.635 1.340 2.050 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.430 0.440 0.670 0.600 ;
    END
END OA31D2

MACRO OA31D4
    CLASS CORE ;
    FOREIGN OA31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.780 1.650 4.110 2.030 ;
        RECT  3.780 0.490 4.110 0.870 ;
        RECT  4.110 0.490 4.530 2.030 ;
        RECT  4.530 1.650 4.690 2.030 ;
        RECT  4.530 0.490 4.690 0.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.480 1.180 1.690 1.340 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.375 2.590 1.515 ;
        RECT  2.590 0.950 2.810 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.970 1.330 1.770 ;
        RECT  1.330 1.650 2.970 1.770 ;
        RECT  2.970 1.005 3.120 1.770 ;
        RECT  3.120 1.180 3.170 1.340 ;
        END
    END A1
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END B
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 0.980 2.820 ;
        RECT  0.980 2.180 1.200 2.820 ;
        RECT  1.200 2.220 2.900 2.820 ;
        RECT  2.900 2.180 3.120 2.820 ;
        RECT  3.120 2.220 3.370 2.820 ;
        RECT  3.370 2.180 3.590 2.820 ;
        RECT  3.590 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.130 0.430 3.370 0.590 ;
        RECT  2.590 0.470 3.130 0.590 ;
        RECT  2.370 0.430 2.590 0.590 ;
        RECT  1.830 0.470 2.370 0.590 ;
        RECT  1.610 0.430 1.830 0.590 ;
        RECT  1.070 0.470 1.610 0.590 ;
        RECT  0.850 0.430 1.070 0.850 ;
        RECT  0.290 0.470 0.850 0.590 ;
        RECT  3.610 1.080 3.890 1.240 ;
        RECT  3.490 0.710 3.610 2.050 ;
        RECT  2.210 0.710 3.490 0.830 ;
        RECT  0.780 1.890 3.490 2.050 ;
        RECT  1.230 0.710 2.210 0.850 ;
        RECT  0.560 1.635 0.780 2.050 ;
        RECT  0.070 0.430 0.290 0.850 ;
        LAYER M1 ;
        RECT  3.780 0.490 3.895 0.870 ;
        RECT  3.780 1.650 3.895 2.030 ;
    END
END OA31D4

MACRO OA32D0
    CLASS CORE ;
    FOREIGN OA32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 0.420 2.470 2.090 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.050 0.640 1.270 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.320 1.050 1.540 ;
        RECT  1.050 1.285 1.190 1.795 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.320 1.370 1.540 ;
        RECT  1.370 1.285 1.510 1.795 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.285 1.830 1.795 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.360 0.300 ;
        RECT  0.360 -0.300 0.580 0.870 ;
        RECT  0.580 -0.300 1.870 0.300 ;
        RECT  1.870 -0.300 2.090 0.340 ;
        RECT  2.090 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.030 0.850 2.190 2.040 ;
        RECT  1.030 0.850 2.030 1.010 ;
        RECT  1.020 1.920 2.030 2.040 ;
        RECT  0.780 1.920 1.020 2.080 ;
    END
END OA32D0

MACRO OA32D1
    CLASS CORE ;
    FOREIGN OA32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 2.200 2.820 ;
        RECT  2.200 2.180 2.420 2.820 ;
        RECT  2.420 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.910 0.440 2.150 0.600 ;
        RECT  1.430 0.480 1.910 0.600 ;
        RECT  1.210 0.440 1.430 0.600 ;
        RECT  0.670 0.480 1.210 0.600 ;
        RECT  2.350 0.720 2.510 1.760 ;
        RECT  0.290 0.720 2.350 0.880 ;
        RECT  1.370 1.640 2.350 1.760 ;
        RECT  1.150 1.640 1.370 2.060 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.430 0.440 0.670 0.600 ;
    END
END OA32D1

MACRO OA32D2
    CLASS CORE ;
    FOREIGN OA32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.560 1.960 2.590 2.100 ;
        RECT  2.590 1.390 2.650 2.100 ;
        RECT  2.590 0.420 2.650 0.900 ;
        RECT  2.650 0.420 2.750 2.100 ;
        RECT  2.750 1.960 2.780 2.100 ;
        RECT  2.750 0.780 2.790 1.515 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.910 0.430 2.150 0.590 ;
        RECT  1.430 0.470 1.910 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  2.310 0.710 2.470 1.760 ;
        RECT  0.290 0.710 2.310 0.870 ;
        RECT  1.370 1.640 2.310 1.760 ;
        RECT  1.150 1.640 1.370 2.060 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  0.430 0.430 0.670 0.590 ;
    END
END OA32D2

MACRO OA32D4
    CLASS CORE ;
    FOREIGN OA32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.390 1.650 4.750 2.030 ;
        RECT  4.390 0.490 4.750 0.870 ;
        RECT  4.750 0.490 5.170 2.030 ;
        RECT  5.170 1.650 5.320 2.030 ;
        RECT  5.170 0.490 5.320 0.870 ;
        END
    END Z
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.260 1.515 ;
        RECT  1.260 1.030 1.420 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.150 2.200 1.515 ;
        RECT  2.200 1.395 3.120 1.515 ;
        RECT  3.120 1.030 3.280 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.800 ;
        RECT  1.850 1.680 3.460 1.800 ;
        RECT  3.460 1.130 3.620 1.800 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 1.440 2.820 ;
        RECT  1.440 2.180 1.660 2.820 ;
        RECT  1.660 2.220 3.590 2.820 ;
        RECT  3.590 2.180 3.810 2.820 ;
        RECT  3.810 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.720 0.430 3.960 0.590 ;
        RECT  3.180 0.470 3.720 0.590 ;
        RECT  2.960 0.430 3.180 0.590 ;
        RECT  2.420 0.470 2.960 0.590 ;
        RECT  2.200 0.430 2.420 0.590 ;
        RECT  1.660 0.470 2.200 0.590 ;
        RECT  1.440 0.430 1.660 0.850 ;
        RECT  0.970 0.470 1.440 0.620 ;
        RECT  0.750 0.430 0.970 0.850 ;
        RECT  0.280 0.470 0.750 0.600 ;
        RECT  4.110 0.710 4.270 2.050 ;
        RECT  1.800 0.710 4.110 0.850 ;
        RECT  2.800 1.930 4.110 2.050 ;
        RECT  2.580 1.930 2.800 2.090 ;
        RECT  0.980 1.930 2.580 2.050 ;
        RECT  0.760 1.635 0.980 2.050 ;
        RECT  0.060 0.420 0.280 0.840 ;
        LAYER M1 ;
        RECT  4.390 0.490 4.535 0.870 ;
        RECT  4.390 1.650 4.535 2.030 ;
    END
END OA32D4

MACRO OA33D0
    CLASS CORE ;
    FOREIGN OA33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.680 2.790 2.030 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.265 1.530 1.795 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.265 1.850 1.795 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.265 2.170 1.795 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.265 1.190 1.795 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.285 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.265 0.250 1.795 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.510 0.300 ;
        RECT  1.510 -0.300 1.730 0.870 ;
        RECT  1.730 -0.300 2.240 0.300 ;
        RECT  2.240 -0.300 2.460 0.340 ;
        RECT  2.460 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 2.170 2.820 ;
        RECT  2.170 2.175 2.390 2.820 ;
        RECT  2.390 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 0.990 2.510 2.040 ;
        RECT  1.010 0.990 2.350 1.110 ;
        RECT  1.360 1.920 2.350 2.040 ;
        RECT  1.120 1.920 1.360 2.080 ;
        RECT  0.070 0.710 0.890 0.870 ;
        RECT  0.890 0.710 1.010 1.110 ;
    END
END OA33D0

MACRO OA33D1
    CLASS CORE ;
    FOREIGN OA33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 1.390 2.660 2.100 ;
        RECT  2.630 0.420 2.660 0.955 ;
        RECT  2.660 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.260 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 2.180 2.820 ;
        RECT  2.180 2.180 2.400 2.820 ;
        RECT  2.400 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.430 2.140 0.590 ;
        RECT  1.430 0.470 1.900 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  2.460 1.050 2.540 1.270 ;
        RECT  2.340 0.710 2.460 1.755 ;
        RECT  0.290 0.710 2.340 0.870 ;
        RECT  1.350 1.635 2.340 1.755 ;
        RECT  1.130 1.635 1.350 2.050 ;
        RECT  0.430 0.430 0.670 0.590 ;
        RECT  0.070 0.450 0.290 0.870 ;
    END
END OA33D1

MACRO OA33D2
    CLASS CORE ;
    FOREIGN OA33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 1.390 2.660 2.100 ;
        RECT  2.630 0.420 2.660 0.955 ;
        RECT  2.660 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.260 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.015 0.300 ;
        RECT  3.015 -0.300 3.235 0.340 ;
        RECT  3.235 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 2.180 2.820 ;
        RECT  2.180 2.180 2.400 2.820 ;
        RECT  2.400 2.220 3.015 2.820 ;
        RECT  3.015 2.180 3.235 2.820 ;
        RECT  3.235 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.430 2.140 0.590 ;
        RECT  1.430 0.470 1.900 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  2.460 1.050 2.540 1.270 ;
        RECT  2.340 0.710 2.460 1.755 ;
        RECT  0.290 0.710 2.340 0.870 ;
        RECT  1.350 1.635 2.340 1.755 ;
        RECT  1.130 1.635 1.350 2.050 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  0.430 0.430 0.670 0.590 ;
    END
END OA33D2

MACRO OA33D4
    CLASS CORE ;
    FOREIGN OA33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.070 1.650 5.390 2.030 ;
        RECT  5.070 0.490 5.390 0.870 ;
        RECT  5.390 0.490 5.810 2.030 ;
        RECT  5.810 1.650 5.980 2.030 ;
        RECT  5.810 0.490 5.980 0.870 ;
        END
    END Z
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 0.970 0.840 1.515 ;
        RECT  0.840 1.380 1.670 1.515 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.130 0.500 1.770 ;
        RECT  0.500 1.650 2.010 1.770 ;
        RECT  2.010 1.005 2.170 1.770 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.180 2.970 1.340 ;
        RECT  2.970 1.005 3.110 1.515 ;
        RECT  3.110 1.395 3.870 1.515 ;
        RECT  3.870 1.030 4.030 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.550 0.970 2.710 1.770 ;
        RECT  2.710 1.650 4.250 1.770 ;
        RECT  4.250 1.005 4.410 1.770 ;
        RECT  4.410 1.005 4.710 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 2.280 2.820 ;
        RECT  2.280 2.180 2.500 2.820 ;
        RECT  2.500 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.430 0.430 4.670 0.590 ;
        RECT  3.890 0.470 4.430 0.590 ;
        RECT  3.670 0.430 3.890 0.590 ;
        RECT  3.130 0.470 3.670 0.590 ;
        RECT  2.910 0.430 3.130 0.590 ;
        RECT  2.370 0.470 2.910 0.590 ;
        RECT  2.150 0.430 2.370 0.850 ;
        RECT  1.680 0.470 2.150 0.630 ;
        RECT  1.460 0.430 1.680 0.850 ;
        RECT  0.970 0.470 1.460 0.630 ;
        RECT  0.750 0.430 0.970 0.850 ;
        RECT  0.280 0.470 0.750 0.630 ;
        RECT  4.950 1.080 5.175 1.240 ;
        RECT  4.830 0.710 4.950 2.050 ;
        RECT  2.530 0.710 4.830 0.850 ;
        RECT  0.060 0.420 0.280 0.840 ;
        RECT  1.110 1.890 4.830 2.050 ;
        LAYER M1 ;
        RECT  5.070 0.490 5.175 0.870 ;
        RECT  5.070 1.650 5.175 2.030 ;
    END
END OA33D4

MACRO OAI211D0
    CLASS CORE ;
    FOREIGN OAI211D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.915 0.590 2.070 ;
        RECT  0.590 1.915 1.310 2.050 ;
        RECT  1.310 1.915 1.370 2.070 ;
        RECT  0.990 0.700 1.370 0.860 ;
        RECT  1.370 0.700 1.530 2.070 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.285 0.550 1.795 ;
        RECT  0.550 1.500 0.740 1.660 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.050 1.250 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 0.870 1.270 ;
        RECT  0.870 1.050 0.930 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.070 0.300 ;
        RECT  0.070 -0.300 0.290 0.340 ;
        RECT  0.290 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.600 2.820 ;
        END
    END VDD
END OAI211D0

MACRO OAI211D1
    CLASS CORE ;
    FOREIGN OAI211D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.650 0.730 2.070 ;
        RECT  0.730 1.650 1.540 1.770 ;
        RECT  1.540 1.650 1.690 2.070 ;
        RECT  1.230 0.720 1.690 0.880 ;
        RECT  1.690 0.720 1.760 2.070 ;
        RECT  1.760 0.720 1.830 1.770 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.890 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.570 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.200 0.300 ;
        RECT  0.200 -0.300 0.420 0.340 ;
        RECT  0.420 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 0.900 2.820 ;
        RECT  0.900 2.180 1.120 2.820 ;
        RECT  1.120 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.630 0.440 1.850 0.600 ;
        RECT  1.090 0.480 1.630 0.600 ;
        RECT  0.870 0.460 1.090 0.880 ;
    END
END OAI211D1

MACRO OAI211D2
    CLASS CORE ;
    FOREIGN OAI211D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.640 0.650 2.060 ;
        RECT  0.650 1.640 1.140 1.760 ;
        RECT  1.140 1.640 1.360 2.060 ;
        RECT  1.360 1.640 2.150 1.760 ;
        RECT  2.150 1.640 2.370 2.060 ;
        RECT  2.370 1.640 2.970 1.760 ;
        RECT  1.750 0.710 2.970 0.870 ;
        RECT  2.970 0.710 3.110 1.760 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.280 1.515 ;
        RECT  1.280 1.030 1.440 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.680 1.005 1.840 1.515 ;
        RECT  1.840 1.395 2.690 1.515 ;
        RECT  2.690 1.030 2.850 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.730 0.300 ;
        RECT  0.730 -0.300 0.950 0.340 ;
        RECT  0.950 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.810 2.820 ;
        RECT  2.810 2.180 3.030 2.820 ;
        RECT  3.030 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.150 0.430 2.370 0.590 ;
        RECT  2.370 0.470 2.910 0.590 ;
        RECT  2.910 0.430 3.130 0.590 ;
        RECT  1.610 0.470 2.150 0.590 ;
        RECT  1.390 0.470 1.610 0.890 ;
        RECT  0.290 0.470 1.390 0.605 ;
        RECT  0.070 0.470 0.290 0.885 ;
    END
END OAI211D2

MACRO OAI211D4
    CLASS CORE ;
    FOREIGN OAI211D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  1.430 1.430 1.870 1.550 ;
        RECT  0.325 0.750 1.870 0.870 ;
        RECT  1.870 0.750 2.290 1.550 ;
        RECT  2.290 0.750 3.365 0.870 ;
        RECT  2.290 1.430 3.790 1.550 ;
        RECT  3.790 1.430 4.010 1.850 ;
        RECT  4.010 1.430 4.480 1.550 ;
        RECT  4.480 1.430 4.700 1.850 ;
        RECT  4.700 1.430 5.280 1.550 ;
        RECT  5.280 1.430 5.500 1.850 ;
        RECT  5.500 1.430 5.970 1.550 ;
        RECT  5.970 1.430 6.190 1.850 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.720 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.390 2.820 ;
        RECT  3.390 2.180 3.610 2.820 ;
        RECT  3.610 2.220 4.880 2.820 ;
        RECT  4.880 2.180 5.100 2.820 ;
        RECT  5.100 2.220 6.370 2.820 ;
        RECT  6.370 2.180 6.590 2.820 ;
        RECT  6.590 2.220 6.720 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.990 1.670 3.210 2.050 ;
        RECT  2.460 1.930 2.990 2.050 ;
        RECT  2.240 1.670 2.460 2.050 ;
        RECT  1.810 1.930 2.240 2.050 ;
        RECT  1.590 1.670 1.810 2.050 ;
        RECT  1.050 1.930 1.590 2.050 ;
        RECT  0.830 1.670 1.050 2.050 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  6.390 0.470 6.610 0.870 ;
        RECT  5.920 0.750 6.390 0.870 ;
        RECT  5.700 0.470 5.920 0.870 ;
        RECT  5.230 0.750 5.700 0.870 ;
        RECT  5.010 0.470 5.230 0.870 ;
        RECT  3.490 0.750 5.010 0.870 ;
        RECT  0.465 0.470 4.870 0.630 ;
        RECT  0.070 1.630 0.290 2.050 ;
        LAYER M1 ;
        RECT  5.970 1.430 6.190 1.850 ;
        RECT  5.500 1.430 5.970 1.550 ;
        RECT  5.280 1.430 5.500 1.850 ;
        RECT  4.700 1.430 5.280 1.550 ;
        RECT  4.480 1.430 4.700 1.850 ;
        RECT  4.010 1.430 4.480 1.550 ;
        RECT  3.790 1.430 4.010 1.850 ;
        RECT  1.430 1.430 1.655 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  0.325 0.750 1.655 0.870 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  2.505 0.750 3.365 0.870 ;
        RECT  2.505 1.430 3.790 1.550 ;
    END
END OAI211D4

MACRO OAI21D0
    CLASS CORE ;
    FOREIGN OAI21D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.890 0.720 2.050 ;
        RECT  0.720 0.660 0.880 2.050 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.550 1.515 ;
        RECT  0.550 1.210 0.580 1.430 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.280 2.820 ;
        END
    END VDD
END OAI21D0

MACRO OAI21D1
    CLASS CORE ;
    FOREIGN OAI21D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.760 ;
        RECT  0.550 0.725 0.730 0.885 ;
        RECT  0.550 1.640 0.790 1.760 ;
        RECT  0.790 1.640 1.010 2.060 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.260 0.300 ;
        RECT  1.260 -0.300 1.480 0.340 ;
        RECT  1.480 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.200 2.820 ;
        RECT  1.200 2.180 1.420 2.820 ;
        RECT  1.420 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.870 0.470 1.090 0.885 ;
        RECT  0.330 0.470 0.870 0.590 ;
        RECT  0.090 0.430 0.330 0.590 ;
    END
END OAI21D1

MACRO OAI21D2
    CLASS CORE ;
    FOREIGN OAI21D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.960 0.500 2.100 ;
        RECT  0.500 1.390 0.660 2.100 ;
        RECT  0.660 1.915 0.690 2.100 ;
        RECT  0.660 1.390 0.730 1.515 ;
        RECT  0.730 0.720 0.870 1.515 ;
        RECT  0.690 1.915 1.520 2.050 ;
        RECT  1.520 1.915 1.760 2.075 ;
        RECT  0.870 0.720 2.130 0.880 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.030 1.200 1.795 ;
        RECT  1.200 1.675 2.010 1.795 ;
        RECT  2.010 1.005 2.150 1.795 ;
        RECT  2.150 1.050 2.190 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.870 2.820 ;
        RECT  0.870 2.180 1.090 2.820 ;
        RECT  1.090 2.220 2.180 2.820 ;
        RECT  2.180 2.180 2.400 2.820 ;
        RECT  2.400 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.270 0.470 2.490 0.890 ;
        RECT  1.730 0.470 2.270 0.590 ;
        RECT  1.510 0.430 1.730 0.590 ;
        RECT  0.970 0.470 1.510 0.590 ;
        RECT  0.750 0.430 0.970 0.590 ;
        RECT  0.280 0.470 0.750 0.590 ;
        RECT  0.060 0.470 0.280 0.885 ;
    END
END OAI21D2

MACRO OAI21D4
    CLASS CORE ;
    FOREIGN OAI21D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  1.430 1.430 1.870 1.550 ;
        RECT  0.325 0.750 1.870 0.870 ;
        RECT  1.870 0.750 2.290 1.550 ;
        RECT  2.290 0.750 3.385 0.870 ;
        RECT  2.290 1.430 3.790 1.550 ;
        RECT  3.790 1.430 4.010 1.850 ;
        RECT  4.010 1.430 4.480 1.550 ;
        RECT  4.480 1.430 4.700 1.850 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END B
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.390 2.820 ;
        RECT  3.390 2.180 3.610 2.820 ;
        RECT  3.610 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.990 1.670 3.210 2.050 ;
        RECT  2.460 1.930 2.990 2.050 ;
        RECT  2.240 1.670 2.460 2.050 ;
        RECT  1.810 1.930 2.240 2.050 ;
        RECT  1.590 1.670 1.810 2.050 ;
        RECT  1.050 1.930 1.590 2.050 ;
        RECT  0.830 1.670 1.050 2.050 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  4.480 0.470 4.700 0.870 ;
        RECT  4.010 0.470 4.480 0.630 ;
        RECT  3.790 0.470 4.010 0.870 ;
        RECT  0.465 0.470 3.790 0.630 ;
        RECT  0.070 1.630 0.290 2.050 ;
        LAYER M1 ;
        RECT  4.480 1.430 4.700 1.850 ;
        RECT  4.010 1.430 4.480 1.550 ;
        RECT  3.790 1.430 4.010 1.850 ;
        RECT  1.430 1.430 1.655 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  0.325 0.750 1.655 0.870 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  2.505 0.750 3.385 0.870 ;
        RECT  2.505 1.430 3.790 1.550 ;
    END
END OAI21D4

MACRO OAI221D0
    CLASS CORE ;
    FOREIGN OAI221D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.910 0.550 2.080 ;
        RECT  0.550 1.920 0.700 2.080 ;
        RECT  0.550 0.910 0.900 1.030 ;
        RECT  0.900 0.710 1.020 1.030 ;
        RECT  1.020 0.710 1.450 0.870 ;
        RECT  0.700 1.920 1.810 2.040 ;
        RECT  1.810 1.920 2.050 2.080 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.490 1.150 1.760 ;
        RECT  1.150 1.640 2.000 1.760 ;
        RECT  2.000 1.005 2.160 1.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.170 1.370 1.390 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.005 1.830 1.515 ;
        END
    END A1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.150 0.870 1.795 ;
        END
    END B2
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.150 2.820 ;
        RECT  1.150 2.180 1.370 2.820 ;
        RECT  1.370 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.690 0.470 1.620 0.590 ;
        RECT  1.620 0.470 1.740 0.820 ;
        RECT  1.740 0.660 2.170 0.820 ;
        RECT  0.470 0.470 0.690 0.790 ;
    END
END OAI221D0

MACRO OAI221D1
    CLASS CORE ;
    FOREIGN OAI221D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.960 0.500 2.100 ;
        RECT  0.500 1.370 0.660 2.100 ;
        RECT  0.660 1.960 0.690 2.100 ;
        RECT  0.660 1.640 1.510 1.760 ;
        RECT  1.510 1.640 1.730 2.060 ;
        RECT  1.730 1.640 2.330 1.760 ;
        RECT  1.880 0.710 2.330 0.870 ;
        RECT  2.330 0.710 2.470 1.760 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.130 2.820 ;
        RECT  1.130 2.180 1.350 2.820 ;
        RECT  1.350 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.180 0.430 1.400 0.590 ;
        RECT  0.640 0.470 1.180 0.590 ;
        RECT  2.280 0.430 2.500 0.590 ;
        RECT  1.740 0.470 2.280 0.590 ;
        RECT  1.520 0.450 1.740 0.870 ;
        RECT  0.420 0.470 0.640 0.885 ;
        RECT  0.780 0.710 1.520 0.870 ;
    END
END OAI221D1

MACRO OAI221D2
    CLASS CORE ;
    FOREIGN OAI221D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  0.100 1.370 0.260 2.100 ;
        RECT  0.260 1.960 0.290 2.100 ;
        RECT  0.260 1.640 0.870 1.760 ;
        RECT  0.870 1.640 1.090 2.060 ;
        RECT  1.090 1.640 2.200 1.760 ;
        RECT  2.200 1.640 2.425 2.060 ;
        RECT  2.425 1.640 2.650 1.760 ;
        RECT  2.650 0.710 2.790 1.760 ;
        RECT  2.790 1.640 3.015 2.060 ;
        RECT  3.015 1.640 4.120 1.760 ;
        RECT  2.790 0.710 4.190 0.870 ;
        RECT  4.120 1.640 4.340 2.060 ;
        RECT  4.190 0.450 4.410 0.870 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.070 1.235 ;
        RECT  1.070 1.005 1.190 1.515 ;
        RECT  1.190 1.395 2.080 1.515 ;
        RECT  2.080 1.030 2.240 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.005 3.110 1.515 ;
        RECT  3.110 1.395 4.000 1.515 ;
        RECT  4.000 1.030 4.160 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.180 0.690 2.820 ;
        RECT  0.690 2.220 1.540 2.820 ;
        RECT  1.540 2.180 1.760 2.820 ;
        RECT  1.760 2.220 3.450 2.820 ;
        RECT  3.450 2.180 3.670 2.820 ;
        RECT  3.670 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.930 0.430 2.150 0.590 ;
        RECT  2.150 0.470 3.050 0.590 ;
        RECT  3.050 0.430 3.270 0.590 ;
        RECT  3.270 0.470 3.810 0.590 ;
        RECT  3.810 0.430 4.050 0.590 ;
        RECT  0.290 0.730 0.790 0.870 ;
        RECT  0.790 0.450 1.010 0.870 ;
        RECT  1.010 0.710 2.530 0.870 ;
        RECT  1.390 0.470 1.930 0.590 ;
        RECT  1.150 0.430 1.390 0.590 ;
        RECT  0.070 0.450 0.290 0.870 ;
    END
END OAI221D2

MACRO OAI221D4
    CLASS CORE ;
    FOREIGN OAI221D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.610 1.640 2.830 2.020 ;
        RECT  2.680 0.760 2.830 0.920 ;
        RECT  2.830 0.760 3.250 2.020 ;
        RECT  3.250 1.640 3.620 2.020 ;
        RECT  3.250 0.760 3.670 0.920 ;
        END
    END ZN
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.240 1.270 ;
        END
    END C
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.160 2.820 ;
        RECT  1.160 2.180 1.380 2.820 ;
        RECT  1.380 2.220 2.220 2.820 ;
        RECT  2.220 2.180 2.440 2.820 ;
        RECT  2.440 2.220 3.000 2.820 ;
        RECT  3.000 2.180 3.220 2.820 ;
        RECT  3.220 2.220 3.790 2.820 ;
        RECT  3.790 2.180 4.010 2.820 ;
        RECT  4.010 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.780 1.635 1.000 2.050 ;
        RECT  1.000 1.635 1.820 1.755 ;
        RECT  1.820 1.635 2.040 2.050 ;
        RECT  2.040 1.635 2.360 1.755 ;
        RECT  2.360 0.470 2.480 1.755 ;
        RECT  2.480 0.470 3.980 0.590 ;
        RECT  3.980 0.470 4.100 1.270 ;
        RECT  4.100 1.050 4.140 1.270 ;
        RECT  1.410 0.470 1.950 0.590 ;
        RECT  1.950 0.470 2.170 0.885 ;
        RECT  0.290 0.470 0.830 0.590 ;
        RECT  0.830 0.470 1.050 0.880 ;
        RECT  1.050 0.720 1.810 0.880 ;
        RECT  0.540 1.635 0.780 1.755 ;
        RECT  0.540 0.720 0.690 0.880 ;
        RECT  4.380 1.960 4.410 2.100 ;
        RECT  4.260 0.420 4.380 2.100 ;
        RECT  4.220 0.420 4.260 0.900 ;
        RECT  4.220 1.390 4.260 2.100 ;
        RECT  3.760 1.390 4.220 1.510 ;
        RECT  4.190 1.960 4.220 2.100 ;
        RECT  3.600 1.050 3.760 1.510 ;
        RECT  0.420 0.720 0.540 1.755 ;
        RECT  1.170 0.430 1.410 0.590 ;
        RECT  0.070 0.470 0.290 0.885 ;
        LAYER M1 ;
        RECT  3.465 1.640 3.620 2.020 ;
        RECT  3.465 0.760 3.670 0.920 ;
        RECT  2.610 1.640 2.615 2.020 ;
    END
END OAI221D4

MACRO OAI222D0
    CLASS CORE ;
    FOREIGN OAI222D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.750 0.870 2.050 ;
        RECT  0.870 0.750 1.530 0.870 ;
        RECT  1.530 0.710 1.770 0.870 ;
        RECT  0.870 1.890 2.360 2.050 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.340 1.490 1.500 1.760 ;
        RECT  1.500 1.640 2.310 1.760 ;
        RECT  2.310 1.005 2.470 1.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.500 1.200 1.690 1.360 ;
        RECT  1.690 1.005 1.830 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.420 0.300 ;
        RECT  0.420 -0.300 0.640 0.340 ;
        RECT  0.640 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.460 2.820 ;
        RECT  1.460 2.180 1.680 2.820 ;
        RECT  1.680 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.260 0.470 0.780 0.590 ;
        RECT  0.780 0.470 1.000 0.630 ;
        RECT  1.000 0.470 2.300 0.590 ;
        RECT  2.300 0.470 2.460 0.870 ;
        RECT  0.100 0.470 0.260 0.870 ;
    END
END OAI222D0

MACRO OAI222D1
    CLASS CORE ;
    FOREIGN OAI222D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.790 1.640 1.010 2.060 ;
        RECT  1.010 1.640 1.850 1.760 ;
        RECT  1.850 1.640 2.070 2.060 ;
        RECT  2.070 1.640 2.330 1.760 ;
        RECT  2.170 0.710 2.330 0.870 ;
        RECT  2.330 0.710 2.470 1.760 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 1.005 1.510 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.005 2.790 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 1.490 2.820 ;
        RECT  1.490 2.180 1.710 2.820 ;
        RECT  1.710 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 2.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.540 0.420 1.780 0.590 ;
        RECT  1.000 0.470 1.540 0.590 ;
        RECT  0.780 0.470 1.000 0.885 ;
        RECT  0.290 0.470 0.780 0.590 ;
        RECT  2.570 0.470 2.810 0.630 ;
        RECT  2.030 0.470 2.570 0.590 ;
        RECT  1.910 0.470 2.030 0.880 ;
        RECT  0.070 0.470 0.290 0.890 ;
        RECT  1.140 0.720 1.910 0.880 ;
    END
END OAI222D1

MACRO OAI222D2
    CLASS CORE ;
    FOREIGN OAI222D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.635 1.020 2.050 ;
        RECT  1.020 1.635 2.200 1.755 ;
        RECT  2.200 1.635 2.420 2.050 ;
        RECT  2.420 1.635 4.060 1.755 ;
        RECT  4.060 1.635 4.280 2.050 ;
        RECT  3.300 0.720 4.840 0.880 ;
        RECT  4.280 1.635 4.870 1.755 ;
        RECT  4.840 0.460 4.870 0.880 ;
        RECT  4.870 0.460 5.030 1.755 ;
        RECT  5.030 0.460 5.060 0.880 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.350 1.515 ;
        RECT  1.350 1.030 1.510 1.515 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.030 1.860 1.515 ;
        RECT  1.860 1.395 2.650 1.515 ;
        RECT  2.650 1.005 2.770 1.515 ;
        RECT  2.770 1.005 3.110 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.590 1.235 ;
        RECT  3.590 1.005 3.750 1.515 ;
        RECT  3.750 1.395 4.570 1.515 ;
        RECT  4.570 1.030 4.730 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.390 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.120 2.820 ;
        RECT  0.120 2.180 0.340 2.820 ;
        RECT  0.340 2.220 1.490 2.820 ;
        RECT  1.490 2.180 1.710 2.820 ;
        RECT  1.710 2.220 2.860 2.820 ;
        RECT  2.860 2.180 3.080 2.820 ;
        RECT  3.080 2.220 3.400 2.820 ;
        RECT  3.400 2.180 3.620 2.820 ;
        RECT  3.620 2.220 4.720 2.820 ;
        RECT  4.720 2.180 4.940 2.820 ;
        RECT  4.940 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.660 0.720 3.180 0.880 ;
        RECT  1.440 0.450 1.660 0.880 ;
        RECT  0.970 0.740 1.440 0.880 ;
        RECT  0.750 0.450 0.970 0.880 ;
        RECT  0.280 0.740 0.750 0.880 ;
        RECT  4.440 0.430 4.680 0.590 ;
        RECT  3.900 0.470 4.440 0.590 ;
        RECT  3.680 0.430 3.900 0.590 ;
        RECT  2.800 0.470 3.680 0.590 ;
        RECT  2.580 0.430 2.800 0.590 ;
        RECT  2.040 0.470 2.580 0.590 ;
        RECT  0.060 0.450 0.280 0.880 ;
        RECT  1.800 0.430 2.040 0.590 ;
    END
END OAI222D2

MACRO OAI222D4
    CLASS CORE ;
    FOREIGN OAI222D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.640 3.150 2.020 ;
        RECT  3.010 0.760 3.150 0.920 ;
        RECT  3.150 0.760 3.570 2.020 ;
        RECT  3.570 1.640 3.950 2.020 ;
        RECT  3.570 0.760 3.990 0.920 ;
        END
    END ZN
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.590 1.270 ;
        END
    END C1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.830 2.820 ;
        RECT  0.830 2.180 1.050 2.820 ;
        RECT  1.050 2.220 2.560 2.820 ;
        RECT  2.560 2.180 2.780 2.820 ;
        RECT  2.780 2.220 3.340 2.820 ;
        RECT  3.340 2.180 3.560 2.820 ;
        RECT  3.560 2.220 4.120 2.820 ;
        RECT  4.120 2.180 4.340 2.820 ;
        RECT  4.340 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.580 0.420 4.700 2.100 ;
        RECT  4.700 1.960 4.730 2.100 ;
        RECT  0.390 1.640 0.450 1.760 ;
        RECT  0.450 0.710 0.570 1.760 ;
        RECT  0.570 0.710 0.690 0.870 ;
        RECT  0.570 1.640 1.500 1.760 ;
        RECT  1.500 1.640 1.720 2.060 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.720 1.640 1.950 1.760 ;
        RECT  1.950 1.370 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 1.640 2.710 1.760 ;
        RECT  2.710 0.470 2.830 1.760 ;
        RECT  2.830 0.470 4.300 0.590 ;
        RECT  4.300 0.470 4.420 1.270 ;
        RECT  4.420 1.050 4.460 1.270 ;
        RECT  2.290 0.460 2.510 0.880 ;
        RECT  0.290 0.470 0.830 0.590 ;
        RECT  0.830 0.470 1.050 0.885 ;
        RECT  1.050 0.470 1.590 0.600 ;
        RECT  1.590 0.440 1.830 0.600 ;
        RECT  4.540 0.420 4.580 0.900 ;
        RECT  4.540 1.390 4.580 2.100 ;
        RECT  4.080 1.390 4.540 1.510 ;
        RECT  4.510 1.960 4.540 2.100 ;
        RECT  3.920 1.050 4.080 1.510 ;
        RECT  0.170 1.640 0.390 2.060 ;
        RECT  1.190 0.720 2.290 0.880 ;
        RECT  0.070 0.470 0.290 0.885 ;
        LAYER M1 ;
        RECT  3.785 1.640 3.950 2.020 ;
        RECT  3.785 0.760 3.990 0.920 ;
    END
END OAI222D4

MACRO OAI22D0
    CLASS CORE ;
    FOREIGN OAI22D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 0.610 0.750 1.235 ;
        RECT  0.750 0.610 0.870 1.810 ;
        RECT  0.870 1.670 0.990 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.510 0.630 2.050 ;
        RECT  0.630 1.930 1.350 2.050 ;
        RECT  1.350 0.790 1.510 2.050 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.570 1.370 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.600 2.820 ;
        END
    END VDD
END OAI22D0

MACRO OAI22D1
    CLASS CORE ;
    FOREIGN OAI22D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.170 1.680 0.390 2.100 ;
        RECT  0.390 1.680 1.510 1.800 ;
        RECT  1.510 1.680 1.690 2.100 ;
        RECT  1.240 0.710 1.690 0.870 ;
        RECT  1.690 0.710 1.730 2.100 ;
        RECT  1.730 0.710 1.830 1.800 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.680 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.350 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.540 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.840 2.820 ;
        RECT  0.840 2.180 1.060 2.820 ;
        RECT  1.060 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.280 0.470 0.880 0.590 ;
        RECT  0.880 0.470 1.100 0.885 ;
        RECT  1.100 0.470 1.640 0.590 ;
        RECT  1.640 0.430 1.860 0.590 ;
        RECT  0.060 0.470 0.280 0.885 ;
    END
END OAI22D1

MACRO OAI22D2
    CLASS CORE ;
    FOREIGN OAI22D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.880 1.640 1.100 2.060 ;
        RECT  1.100 1.640 1.690 1.760 ;
        RECT  1.690 0.720 1.830 1.760 ;
        RECT  1.830 1.640 2.440 1.760 ;
        RECT  2.440 1.640 2.660 2.060 ;
        RECT  1.830 0.720 3.060 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        RECT  0.560 1.395 1.410 1.515 ;
        RECT  1.410 1.030 1.570 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.950 1.030 2.110 1.515 ;
        RECT  2.110 1.395 2.960 1.515 ;
        RECT  2.960 1.005 3.120 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.790 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.700 0.340 ;
        RECT  0.700 -0.300 1.280 0.300 ;
        RECT  1.280 -0.300 1.500 0.340 ;
        RECT  1.500 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.220 2.820 ;
        RECT  0.220 2.180 0.440 2.820 ;
        RECT  0.440 2.220 1.670 2.820 ;
        RECT  1.670 2.180 1.890 2.820 ;
        RECT  1.890 2.220 3.100 2.820 ;
        RECT  3.100 2.180 3.320 2.820 ;
        RECT  3.320 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.200 0.470 3.420 0.890 ;
        RECT  2.660 0.470 3.200 0.590 ;
        RECT  2.440 0.430 2.660 0.590 ;
        RECT  1.900 0.470 2.440 0.590 ;
        RECT  1.680 0.430 1.900 0.590 ;
        RECT  1.100 0.470 1.680 0.590 ;
        RECT  0.880 0.470 1.100 0.885 ;
        RECT  0.300 0.470 0.880 0.590 ;
        RECT  0.080 0.470 0.300 0.890 ;
    END
END OAI22D2

MACRO OAI22D4
    CLASS CORE ;
    FOREIGN OAI22D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  1.430 1.430 1.870 1.550 ;
        RECT  0.325 0.750 1.870 0.870 ;
        RECT  1.870 0.750 2.290 1.550 ;
        RECT  2.290 0.750 3.385 0.870 ;
        RECT  2.290 1.430 5.580 1.550 ;
        RECT  5.580 1.430 5.800 1.810 ;
        RECT  5.800 1.430 6.340 1.550 ;
        RECT  6.340 1.430 6.560 1.810 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.710 1.235 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 6.310 1.235 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.505 0.300 ;
        RECT  3.505 -0.300 3.725 0.340 ;
        RECT  3.725 -0.300 4.300 0.300 ;
        RECT  4.300 -0.300 4.520 0.340 ;
        RECT  4.520 -0.300 5.090 0.300 ;
        RECT  5.090 -0.300 5.310 0.340 ;
        RECT  5.310 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.340 ;
        RECT  6.110 -0.300 6.690 0.300 ;
        RECT  6.690 -0.300 6.910 0.340 ;
        RECT  6.910 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 3.400 2.820 ;
        RECT  3.400 2.180 3.620 2.820 ;
        RECT  3.620 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.000 1.670 3.220 2.050 ;
        RECT  2.460 1.930 3.000 2.050 ;
        RECT  2.240 1.670 2.460 2.050 ;
        RECT  1.810 1.930 2.240 2.050 ;
        RECT  1.590 1.670 1.810 2.050 ;
        RECT  1.050 1.930 1.590 2.050 ;
        RECT  0.830 1.670 1.050 2.050 ;
        RECT  0.290 1.930 0.830 2.050 ;
        RECT  6.290 0.470 6.510 0.870 ;
        RECT  5.710 0.470 6.290 0.630 ;
        RECT  5.490 0.470 5.710 0.870 ;
        RECT  4.910 0.470 5.490 0.630 ;
        RECT  4.690 0.470 4.910 0.870 ;
        RECT  4.125 0.470 4.690 0.630 ;
        RECT  3.905 0.470 4.125 0.870 ;
        RECT  6.720 1.630 6.940 2.050 ;
        RECT  6.180 1.930 6.720 2.050 ;
        RECT  5.960 1.670 6.180 2.050 ;
        RECT  5.420 1.930 5.960 2.050 ;
        RECT  5.200 1.670 5.420 2.050 ;
        RECT  4.780 1.930 5.200 2.050 ;
        RECT  4.560 1.670 4.780 2.050 ;
        RECT  4.020 1.930 4.560 2.050 ;
        RECT  0.465 0.470 3.905 0.630 ;
        RECT  0.070 1.630 0.290 2.050 ;
        RECT  3.800 1.670 4.020 2.050 ;
        LAYER M1 ;
        RECT  6.340 1.430 6.560 1.810 ;
        RECT  5.800 1.430 6.340 1.550 ;
        RECT  5.580 1.430 5.800 1.810 ;
        RECT  1.430 1.430 1.655 1.550 ;
        RECT  1.210 1.430 1.430 1.810 ;
        RECT  0.670 1.430 1.210 1.550 ;
        RECT  0.325 0.750 1.655 0.870 ;
        RECT  0.105 0.470 0.325 0.870 ;
        RECT  0.450 1.430 0.670 1.810 ;
        RECT  2.505 0.750 3.385 0.870 ;
        RECT  2.505 1.430 5.580 1.550 ;
    END
END OAI22D4

MACRO OAI31D0
    CLASS CORE ;
    FOREIGN OAI31D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.490 0.260 0.880 ;
        RECT  0.260 0.760 0.840 0.880 ;
        RECT  0.840 0.710 1.060 0.880 ;
        RECT  1.110 1.860 1.690 2.020 ;
        RECT  1.060 0.760 1.690 0.880 ;
        RECT  1.690 0.760 1.830 2.020 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.540 2.820 ;
        RECT  1.540 2.180 1.760 2.820 ;
        RECT  1.760 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.230 0.470 1.470 0.640 ;
        RECT  0.670 0.470 1.230 0.590 ;
        RECT  0.430 0.470 0.670 0.640 ;
    END
END OAI31D0

MACRO OAI31D1
    CLASS CORE ;
    FOREIGN OAI31D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  1.130 1.640 1.350 2.060 ;
        RECT  1.350 1.640 1.690 1.760 ;
        RECT  0.290 0.710 1.690 0.870 ;
        RECT  1.690 0.710 1.830 1.760 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.510 1.515 ;
        RECT  1.510 1.050 1.530 1.270 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.160 2.820 ;
        RECT  0.160 2.180 0.380 2.820 ;
        RECT  0.380 2.220 1.540 2.820 ;
        RECT  1.540 2.180 1.760 2.820 ;
        RECT  1.760 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.210 0.430 1.450 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  0.430 0.430 0.670 0.590 ;
    END
END OAI31D1

MACRO OAI31D2
    CLASS CORE ;
    FOREIGN OAI31D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.630 0.860 2.050 ;
        RECT  0.860 1.890 3.290 2.050 ;
        RECT  1.310 0.710 3.290 0.860 ;
        RECT  3.290 0.710 3.430 2.050 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.570 1.515 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.630 1.140 1.790 1.515 ;
        RECT  1.790 1.395 2.650 1.515 ;
        RECT  2.650 1.005 2.810 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.390 1.235 ;
        RECT  1.390 1.005 1.510 1.760 ;
        RECT  1.510 1.640 3.010 1.760 ;
        RECT  3.010 1.140 3.170 1.760 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.530 0.300 ;
        RECT  0.530 -0.300 0.750 0.340 ;
        RECT  0.750 -0.300 3.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.230 2.820 ;
        RECT  0.230 2.180 0.450 2.820 ;
        RECT  0.450 2.220 1.050 2.820 ;
        RECT  1.050 2.180 1.270 2.820 ;
        RECT  1.270 2.220 3.150 2.820 ;
        RECT  3.150 2.180 3.370 2.820 ;
        RECT  3.370 2.220 3.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.230 0.430 3.450 0.590 ;
        RECT  2.690 0.470 3.230 0.590 ;
        RECT  2.470 0.430 2.690 0.590 ;
        RECT  1.930 0.470 2.470 0.590 ;
        RECT  1.710 0.430 1.930 0.590 ;
        RECT  1.170 0.470 1.710 0.590 ;
        RECT  0.950 0.440 1.170 0.860 ;
        RECT  0.340 0.470 0.950 0.600 ;
        RECT  0.120 0.440 0.340 0.860 ;
    END
END OAI31D2

MACRO OAI31D4
    CLASS CORE ;
    FOREIGN OAI31D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.040 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.145 0.470 0.365 0.870 ;
        RECT  0.490 1.430 0.710 1.810 ;
        RECT  0.710 1.430 1.250 1.550 ;
        RECT  1.250 1.430 1.470 1.810 ;
        RECT  1.470 1.430 3.790 1.550 ;
        RECT  0.365 0.750 3.790 0.870 ;
        RECT  3.790 0.750 4.210 1.550 ;
        RECT  4.210 0.750 5.305 0.870 ;
        RECT  4.210 1.430 5.710 1.550 ;
        RECT  5.710 1.430 5.930 1.850 ;
        RECT  5.930 1.430 6.400 1.550 ;
        RECT  6.400 1.430 6.620 1.850 ;
        END
    END ZN
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.005 6.630 1.235 ;
        END
    END B
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 7.040 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.310 2.820 ;
        RECT  5.310 2.180 5.530 2.820 ;
        RECT  5.530 2.220 7.040 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.850 1.670 3.370 1.810 ;
        RECT  1.630 1.670 1.850 2.050 ;
        RECT  1.090 1.930 1.630 2.050 ;
        RECT  0.870 1.670 1.090 2.050 ;
        RECT  0.330 1.930 0.870 2.050 ;
        RECT  4.910 1.670 5.130 2.050 ;
        RECT  4.380 1.930 4.910 2.050 ;
        RECT  4.160 1.670 4.380 2.050 ;
        RECT  3.730 1.930 4.160 2.050 ;
        RECT  3.510 1.670 3.730 2.050 ;
        RECT  6.400 0.470 6.620 0.870 ;
        RECT  5.930 0.470 6.400 0.630 ;
        RECT  5.710 0.470 5.930 0.870 ;
        RECT  0.505 0.470 5.710 0.630 ;
        RECT  1.970 1.930 3.510 2.050 ;
        RECT  0.110 1.630 0.330 2.050 ;
        LAYER M1 ;
        RECT  6.400 1.430 6.620 1.850 ;
        RECT  5.930 1.430 6.400 1.550 ;
        RECT  5.710 1.430 5.930 1.850 ;
        RECT  1.470 1.430 3.575 1.550 ;
        RECT  1.250 1.430 1.470 1.810 ;
        RECT  0.710 1.430 1.250 1.550 ;
        RECT  0.365 0.750 3.575 0.870 ;
        RECT  0.145 0.470 0.365 0.870 ;
        RECT  0.490 1.430 0.710 1.810 ;
        RECT  4.425 0.750 5.305 0.870 ;
        RECT  4.425 1.430 5.710 1.550 ;
    END
END OAI31D4

MACRO OAI32D0
    CLASS CORE ;
    FOREIGN OAI32D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.440 0.260 0.850 ;
        RECT  1.190 1.880 2.010 2.040 ;
        RECT  0.260 0.710 2.010 0.850 ;
        RECT  2.010 0.710 2.150 2.040 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.250 1.890 1.470 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 1.880 2.820 ;
        RECT  1.880 2.180 2.100 2.820 ;
        RECT  2.100 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.950 0.450 2.170 0.590 ;
        RECT  1.450 0.470 1.950 0.590 ;
        RECT  1.230 0.450 1.450 0.590 ;
        RECT  0.670 0.470 1.230 0.590 ;
        RECT  0.430 0.450 0.670 0.590 ;
    END
END OAI32D0

MACRO OAI32D1
    CLASS CORE ;
    FOREIGN OAI32D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  1.150 1.635 1.370 2.050 ;
        RECT  1.370 1.635 2.010 1.755 ;
        RECT  0.290 0.710 2.010 0.870 ;
        RECT  2.010 0.710 2.150 1.755 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.890 1.270 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 1.860 2.820 ;
        RECT  1.860 2.180 2.080 2.820 ;
        RECT  2.080 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.930 0.430 2.170 0.590 ;
        RECT  1.430 0.470 1.930 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  0.430 0.430 0.670 0.590 ;
    END
END OAI32D1

MACRO OAI32D2
    CLASS CORE ;
    FOREIGN OAI32D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.635 1.050 2.050 ;
        RECT  1.050 1.890 3.930 2.050 ;
        RECT  1.950 0.710 3.930 0.860 ;
        RECT  3.930 0.710 4.070 2.050 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 1.190 1.235 ;
        END
    END B2
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.005 3.110 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.160 2.330 1.380 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.395 3.290 1.515 ;
        RECT  3.290 1.030 3.450 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.030 1.235 ;
        RECT  2.030 1.005 2.150 1.760 ;
        RECT  2.150 1.640 3.610 1.760 ;
        RECT  3.610 1.160 3.750 1.760 ;
        RECT  3.750 1.160 3.810 1.380 ;
        END
    END A1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        RECT  0.550 1.380 1.340 1.515 ;
        RECT  1.340 1.060 1.500 1.515 ;
        END
    END B1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.170 2.820 ;
        RECT  0.170 2.180 0.390 2.820 ;
        RECT  0.390 2.220 1.620 2.820 ;
        RECT  1.620 2.180 1.840 2.820 ;
        RECT  1.840 2.220 3.800 2.820 ;
        RECT  3.800 2.180 4.020 2.820 ;
        RECT  4.020 2.220 4.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.830 0.440 1.050 0.860 ;
        RECT  1.050 0.470 1.590 0.600 ;
        RECT  1.590 0.440 1.810 0.860 ;
        RECT  1.810 0.470 2.350 0.590 ;
        RECT  2.350 0.430 2.570 0.590 ;
        RECT  2.570 0.470 3.110 0.590 ;
        RECT  3.110 0.430 3.330 0.590 ;
        RECT  3.330 0.470 3.870 0.590 ;
        RECT  3.870 0.430 4.090 0.590 ;
        RECT  0.290 0.470 0.830 0.600 ;
        RECT  0.070 0.440 0.290 0.860 ;
    END
END OAI32D2

MACRO OAI32D4
    CLASS CORE ;
    FOREIGN OAI32D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.640 3.470 2.020 ;
        RECT  2.970 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 3.970 2.020 ;
        RECT  3.890 0.500 3.970 0.880 ;
        END
    END ZN
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.580 0.300 ;
        RECT  2.580 -0.300 2.800 0.340 ;
        RECT  2.800 -0.300 3.360 0.300 ;
        RECT  3.360 -0.300 3.580 0.340 ;
        RECT  3.580 -0.300 4.140 0.300 ;
        RECT  4.140 -0.300 4.360 0.340 ;
        RECT  4.360 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 1.850 2.820 ;
        RECT  1.850 2.180 2.070 2.820 ;
        RECT  2.070 2.220 2.580 2.820 ;
        RECT  2.580 2.180 2.800 2.820 ;
        RECT  2.800 2.220 3.360 2.820 ;
        RECT  3.360 2.180 3.580 2.820 ;
        RECT  3.580 2.220 4.140 2.820 ;
        RECT  4.140 2.180 4.360 2.820 ;
        RECT  4.360 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.900 0.430 2.140 0.590 ;
        RECT  1.430 0.470 1.900 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  2.090 1.080 2.560 1.240 ;
        RECT  1.970 0.710 2.090 1.765 ;
        RECT  0.290 0.710 1.970 0.870 ;
        RECT  1.365 1.635 1.970 1.765 ;
        RECT  1.145 1.635 1.365 2.050 ;
        RECT  2.800 1.080 3.080 1.240 ;
        RECT  2.680 0.730 2.800 1.510 ;
        RECT  2.220 0.730 2.680 0.950 ;
        RECT  2.380 1.390 2.680 1.510 ;
        RECT  2.380 1.960 2.410 2.100 ;
        RECT  2.220 1.390 2.380 2.100 ;
        RECT  0.070 0.420 0.290 0.870 ;
        RECT  0.430 0.430 0.670 0.590 ;
        RECT  2.190 1.960 2.220 2.100 ;
        LAYER M1 ;
        RECT  2.970 0.500 3.255 0.880 ;
        RECT  2.970 1.640 3.255 2.020 ;
    END
END OAI32D4

MACRO OAI33D0
    CLASS CORE ;
    FOREIGN OAI33D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.100 0.490 0.260 0.870 ;
        RECT  0.260 0.750 0.840 0.870 ;
        RECT  0.840 0.710 1.060 0.870 ;
        RECT  1.150 1.820 2.330 1.980 ;
        RECT  1.060 0.750 2.330 0.870 ;
        RECT  2.330 0.750 2.470 1.980 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 0.995 1.530 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.850 1.535 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.295 2.200 1.515 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.535 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.535 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.535 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 0.470 2.160 0.630 ;
        RECT  1.450 0.470 1.920 0.590 ;
        RECT  1.230 0.470 1.450 0.630 ;
        RECT  0.670 0.470 1.230 0.590 ;
        RECT  0.430 0.470 0.670 0.630 ;
    END
END OAI33D0

MACRO OAI33D1
    CLASS CORE ;
    FOREIGN OAI33D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.070 0.450 0.290 0.870 ;
        RECT  1.130 1.635 1.350 2.050 ;
        RECT  1.350 1.635 2.330 1.755 ;
        RECT  0.290 0.710 2.330 0.870 ;
        RECT  2.330 0.710 2.470 1.755 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.870 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.050 2.200 1.270 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.370 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.920 0.430 2.160 0.590 ;
        RECT  1.430 0.470 1.920 0.590 ;
        RECT  1.210 0.430 1.430 0.590 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  0.430 0.430 0.670 0.590 ;
    END
END OAI33D1

MACRO OAI33D2
    CLASS CORE ;
    FOREIGN OAI33D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.890 4.570 2.050 ;
        RECT  2.590 0.710 4.570 0.860 ;
        RECT  4.570 0.710 4.710 2.050 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.750 1.235 ;
        RECT  0.750 1.005 0.870 1.475 ;
        RECT  0.870 1.355 1.680 1.475 ;
        RECT  1.680 1.140 1.840 1.475 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.720 ;
        RECT  0.250 1.600 2.030 1.720 ;
        RECT  2.030 0.995 2.190 1.720 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.750 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.160 2.970 1.380 ;
        RECT  2.970 1.005 3.110 1.515 ;
        RECT  3.110 1.395 3.930 1.515 ;
        RECT  3.930 1.030 4.090 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.670 1.235 ;
        RECT  2.670 1.005 2.790 1.760 ;
        RECT  2.790 1.640 4.290 1.760 ;
        RECT  4.290 1.140 4.450 1.760 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.140 2.820 ;
        RECT  0.140 2.180 0.360 2.820 ;
        RECT  0.360 2.220 2.250 2.820 ;
        RECT  2.250 2.180 2.470 2.820 ;
        RECT  2.470 2.220 4.430 2.820 ;
        RECT  4.430 2.180 4.650 2.820 ;
        RECT  4.650 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.290 0.470 0.790 0.600 ;
        RECT  0.790 0.440 1.010 0.860 ;
        RECT  1.010 0.470 1.510 0.600 ;
        RECT  1.510 0.440 1.730 0.860 ;
        RECT  1.730 0.470 2.230 0.600 ;
        RECT  2.230 0.440 2.450 0.860 ;
        RECT  2.450 0.470 2.990 0.590 ;
        RECT  2.990 0.430 3.210 0.590 ;
        RECT  3.210 0.470 3.750 0.590 ;
        RECT  3.750 0.430 3.970 0.590 ;
        RECT  3.970 0.470 4.510 0.590 ;
        RECT  4.510 0.430 4.730 0.590 ;
        RECT  0.070 0.440 0.290 0.860 ;
    END
END OAI33D2

MACRO OAI33D4
    CLASS CORE ;
    FOREIGN OAI33D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 1.640 2.830 2.020 ;
        RECT  2.610 0.760 2.830 0.920 ;
        RECT  2.830 0.760 3.250 2.020 ;
        RECT  3.250 1.640 3.630 2.020 ;
        RECT  3.250 0.760 3.630 0.920 ;
        END
    END ZN
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.530 1.515 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.880 1.270 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.150 1.515 ;
        RECT  2.150 1.080 2.250 1.240 ;
        END
    END B1
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.005 1.200 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.020 0.300 ;
        RECT  3.020 -0.300 3.240 0.340 ;
        RECT  3.240 -0.300 3.800 0.300 ;
        RECT  3.800 -0.300 4.020 0.340 ;
        RECT  4.020 -0.300 4.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.180 2.820 ;
        RECT  0.180 2.180 0.400 2.820 ;
        RECT  0.400 2.220 2.220 2.820 ;
        RECT  2.220 2.180 2.440 2.820 ;
        RECT  2.440 2.220 3.020 2.820 ;
        RECT  3.020 2.180 3.240 2.820 ;
        RECT  3.240 2.220 3.800 2.820 ;
        RECT  3.800 2.180 4.020 2.820 ;
        RECT  4.020 2.220 4.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.540 1.635 1.180 1.755 ;
        RECT  1.180 1.635 1.400 2.050 ;
        RECT  1.400 1.635 2.370 1.755 ;
        RECT  2.370 0.470 2.490 1.755 ;
        RECT  2.490 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.100 1.270 ;
        RECT  0.670 0.470 1.210 0.590 ;
        RECT  1.210 0.470 1.430 0.885 ;
        RECT  1.430 0.470 1.930 0.590 ;
        RECT  1.930 0.470 2.150 0.885 ;
        RECT  0.540 0.720 1.070 0.880 ;
        RECT  0.420 0.720 0.540 1.755 ;
        RECT  0.290 0.720 0.420 0.880 ;
        RECT  4.380 1.960 4.410 2.100 ;
        RECT  4.220 0.420 4.380 2.100 ;
        RECT  3.750 1.390 4.220 1.510 ;
        RECT  4.190 1.960 4.220 2.100 ;
        RECT  3.590 1.050 3.750 1.510 ;
        RECT  0.070 0.460 0.290 0.880 ;
        RECT  0.430 0.430 0.670 0.590 ;
        LAYER M1 ;
        RECT  3.465 1.640 3.630 2.020 ;
        RECT  3.465 0.760 3.630 0.920 ;
    END
END OAI33D4

MACRO OR2D0
    CLASS CORE ;
    FOREIGN OR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.350 0.450 1.510 2.080 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.900 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.920 0.300 ;
        RECT  0.920 -0.300 1.140 0.340 ;
        RECT  1.140 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.910 2.820 ;
        RECT  0.910 2.180 1.130 2.820 ;
        RECT  1.130 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.220 1.870 1.070 2.030 ;
        RECT  0.500 0.540 1.070 0.700 ;
        RECT  1.070 0.540 1.230 2.030 ;
    END
END OR2D0

MACRO OR2D1
    CLASS CORE ;
    FOREIGN OR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.960 1.350 2.100 ;
        RECT  1.350 0.420 1.510 2.100 ;
        RECT  1.510 1.960 1.540 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.900 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.910 0.300 ;
        RECT  0.910 -0.300 1.130 0.340 ;
        RECT  1.130 -0.300 1.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.910 2.820 ;
        RECT  0.910 2.180 1.130 2.820 ;
        RECT  1.130 2.220 1.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.240 1.640 0.460 2.060 ;
        RECT  0.460 1.640 1.070 1.800 ;
        RECT  0.470 0.710 1.070 0.870 ;
        RECT  1.070 0.710 1.230 1.800 ;
    END
END OR2D1

MACRO OR2D2
    CLASS CORE ;
    FOREIGN OR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.280 1.960 1.310 2.100 ;
        RECT  1.310 1.390 1.370 2.100 ;
        RECT  1.310 0.420 1.370 0.900 ;
        RECT  1.370 0.420 1.470 2.100 ;
        RECT  1.470 1.960 1.500 2.100 ;
        RECT  1.470 0.780 1.510 1.515 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.890 0.300 ;
        RECT  0.890 -0.300 1.110 0.340 ;
        RECT  1.110 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.870 2.820 ;
        RECT  0.870 2.180 1.090 2.820 ;
        RECT  1.090 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.030 0.710 1.190 1.760 ;
        RECT  0.470 0.710 1.030 0.870 ;
        RECT  0.420 1.640 1.030 1.760 ;
        RECT  0.200 1.640 0.420 2.060 ;
    END
END OR2D2

MACRO OR2D4
    CLASS CORE ;
    FOREIGN OR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.650 2.190 2.030 ;
        RECT  1.810 0.490 2.190 0.870 ;
        RECT  2.190 0.490 2.610 2.030 ;
        RECT  2.610 1.650 2.720 2.030 ;
        RECT  2.610 0.490 2.720 0.870 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        RECT  0.250 1.395 1.280 1.515 ;
        RECT  1.280 1.030 1.440 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.870 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.770 0.300 ;
        RECT  0.770 -0.300 0.990 0.340 ;
        RECT  0.990 -0.300 1.410 0.300 ;
        RECT  1.410 -0.300 1.630 0.340 ;
        RECT  1.630 -0.300 3.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.130 2.820 ;
        RECT  0.130 2.180 0.350 2.820 ;
        RECT  0.350 2.220 1.420 2.820 ;
        RECT  1.420 2.180 1.640 2.820 ;
        RECT  1.640 2.220 3.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.690 1.080 1.920 1.240 ;
        RECT  1.570 0.710 1.690 1.800 ;
        RECT  0.400 0.710 1.570 0.870 ;
        RECT  0.990 1.640 1.570 1.800 ;
        RECT  0.770 1.640 0.990 2.060 ;
        LAYER M1 ;
        RECT  1.810 0.490 1.975 0.870 ;
        RECT  1.810 1.650 1.975 2.030 ;
    END
END OR2D4

MACRO OR2D8
    CLASS CORE ;
    FOREIGN OR2D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.120 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.640 3.470 2.020 ;
        RECT  2.380 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 4.670 2.020 ;
        RECT  3.890 0.500 4.670 0.880 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.100 0.890 1.800 ;
        RECT  0.890 1.395 1.860 1.515 ;
        RECT  1.860 1.030 2.020 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 0.860 0.460 1.350 ;
        RECT  0.460 0.860 1.050 0.980 ;
        RECT  1.050 0.860 1.170 1.235 ;
        RECT  1.170 1.005 1.510 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.575 0.300 ;
        RECT  0.575 -0.300 0.795 0.340 ;
        RECT  0.795 -0.300 5.120 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.990 2.820 ;
        RECT  1.990 2.180 2.210 2.820 ;
        RECT  2.210 2.220 5.120 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.260 1.080 3.060 1.240 ;
        RECT  2.140 0.520 2.260 2.050 ;
        RECT  0.950 0.520 2.140 0.680 ;
        RECT  1.570 1.930 2.140 2.050 ;
        RECT  1.350 1.650 1.570 2.050 ;
        RECT  0.340 1.930 1.350 2.050 ;
        RECT  0.120 1.650 0.340 2.050 ;
        LAYER M1 ;
        RECT  2.380 0.500 3.255 0.880 ;
        RECT  2.380 1.640 3.255 2.020 ;
        RECT  4.105 0.500 4.670 0.880 ;
        RECT  4.105 1.640 4.670 2.020 ;
    END
END OR2D8

MACRO OR3D0
    CLASS CORE ;
    FOREIGN OR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.600 1.830 1.990 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.250 1.220 1.470 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.230 2.820 ;
        RECT  1.230 2.180 1.450 2.820 ;
        RECT  1.450 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.700 1.550 1.940 ;
        RECT  0.070 0.700 1.390 0.860 ;
        RECT  0.290 1.780 1.390 1.940 ;
    END
END OR3D0

MACRO OR3D1
    CLASS CORE ;
    FOREIGN OR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.640 1.960 1.670 2.100 ;
        RECT  1.670 0.420 1.830 2.100 ;
        RECT  1.830 1.960 1.860 2.100 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.900 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.050 1.220 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 1.250 0.300 ;
        RECT  1.250 -0.300 1.470 0.340 ;
        RECT  1.470 -0.300 1.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.230 2.820 ;
        RECT  1.230 2.180 1.450 2.820 ;
        RECT  1.450 2.220 1.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.390 0.710 1.550 1.760 ;
        RECT  0.070 0.710 1.390 0.870 ;
        RECT  0.460 1.640 1.390 1.760 ;
        RECT  0.240 1.640 0.460 2.060 ;
    END
END OR3D1

MACRO OR3D2
    CLASS CORE ;
    FOREIGN OR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.960 1.630 2.100 ;
        RECT  1.630 1.390 1.690 2.100 ;
        RECT  1.630 0.420 1.690 0.900 ;
        RECT  1.690 0.420 1.790 2.100 ;
        RECT  1.790 1.960 1.820 2.100 ;
        RECT  1.790 0.780 1.830 1.515 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.005 0.870 1.515 ;
        RECT  0.870 1.050 0.900 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.190 1.515 ;
        RECT  1.190 1.050 1.220 1.270 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.340 ;
        RECT  0.680 -0.300 1.200 0.300 ;
        RECT  1.200 -0.300 1.420 0.340 ;
        RECT  1.420 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.210 2.820 ;
        RECT  1.210 2.180 1.430 2.820 ;
        RECT  1.430 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.510 1.050 1.550 1.270 ;
        RECT  1.390 0.710 1.510 1.760 ;
        RECT  0.070 0.710 1.390 0.870 ;
        RECT  0.460 1.640 1.390 1.760 ;
        RECT  0.240 1.640 0.460 2.060 ;
    END
END OR3D2

MACRO OR3D4
    CLASS CORE ;
    FOREIGN OR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.500 1.650 2.830 2.030 ;
        RECT  2.500 0.490 2.830 0.870 ;
        RECT  2.830 0.490 3.250 2.030 ;
        RECT  3.250 1.650 3.410 2.030 ;
        RECT  3.250 0.490 3.410 0.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.005 0.750 1.235 ;
        RECT  0.750 0.765 0.870 1.235 ;
        RECT  0.870 0.765 1.570 0.885 ;
        RECT  1.570 0.765 1.690 1.240 ;
        RECT  1.690 1.080 1.830 1.240 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.755 ;
        RECT  0.250 1.635 1.950 1.755 ;
        RECT  1.950 1.030 2.110 1.755 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.150 2.820 ;
        RECT  0.150 2.180 0.370 2.820 ;
        RECT  0.370 2.220 2.090 2.820 ;
        RECT  2.090 2.180 2.310 2.820 ;
        RECT  2.310 2.220 3.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.350 1.080 2.610 1.240 ;
        RECT  2.230 0.470 2.350 2.050 ;
        RECT  0.410 0.470 2.230 0.630 ;
        RECT  1.100 1.890 2.230 2.050 ;
        LAYER M1 ;
        RECT  2.500 0.490 2.615 0.870 ;
        RECT  2.500 1.650 2.615 2.030 ;
    END
END OR3D4

MACRO OR3D8
    CLASS CORE ;
    FOREIGN OR3D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.480 1.640 4.430 2.020 ;
        RECT  3.540 0.500 4.430 0.880 ;
        RECT  4.430 0.500 4.850 2.020 ;
        RECT  4.850 1.640 5.980 2.020 ;
        RECT  4.850 0.500 5.980 0.880 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.090 0.870 1.250 ;
        RECT  0.870 0.970 0.990 1.250 ;
        RECT  0.990 0.970 1.460 1.090 ;
        RECT  1.460 0.970 1.580 1.125 ;
        RECT  1.580 1.005 1.690 1.125 ;
        RECT  1.690 1.005 2.160 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.510 0.725 0.750 0.870 ;
        RECT  0.750 0.725 1.680 0.845 ;
        RECT  1.680 0.725 2.620 0.870 ;
        RECT  2.620 0.725 2.650 0.890 ;
        RECT  2.650 0.725 2.790 1.235 ;
        RECT  2.790 0.725 2.840 0.890 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.210 1.190 1.350 ;
        RECT  1.190 1.210 1.330 1.680 ;
        RECT  1.330 1.560 2.960 1.680 ;
        RECT  2.960 1.005 3.120 1.680 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.100 2.820 ;
        RECT  1.100 2.180 1.320 2.820 ;
        RECT  1.320 2.220 3.070 2.820 ;
        RECT  3.070 2.180 3.290 2.820 ;
        RECT  3.290 2.220 6.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.360 1.060 4.175 1.220 ;
        RECT  3.240 0.470 3.360 2.050 ;
        RECT  0.060 0.470 3.240 0.590 ;
        RECT  0.360 1.890 3.240 2.050 ;
        RECT  0.140 1.630 0.360 2.050 ;
        LAYER M1 ;
        RECT  3.480 1.640 4.215 2.020 ;
        RECT  3.540 0.500 4.215 0.880 ;
        RECT  5.065 0.500 5.980 0.880 ;
        RECT  5.065 1.640 5.980 2.020 ;
    END
END OR3D8

MACRO OR4D0
    CLASS CORE ;
    FOREIGN OR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.990 0.620 2.150 1.850 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.795 0.300 ;
        RECT  0.795 -0.300 1.015 0.340 ;
        RECT  1.015 -0.300 1.550 0.300 ;
        RECT  1.550 -0.300 1.770 0.340 ;
        RECT  1.770 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.520 2.820 ;
        RECT  1.520 2.180 1.740 2.820 ;
        RECT  1.740 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.710 0.720 1.870 1.800 ;
        RECT  0.190 1.640 1.710 1.800 ;
        RECT  0.430 0.720 1.710 0.880 ;
    END
END OR4D0

MACRO OR4D1
    CLASS CORE ;
    FOREIGN OR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.960 1.990 2.100 ;
        RECT  1.990 0.420 2.150 2.100 ;
        RECT  2.150 1.960 2.180 2.100 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.795 0.300 ;
        RECT  0.795 -0.300 1.015 0.340 ;
        RECT  1.015 -0.300 1.550 0.300 ;
        RECT  1.550 -0.300 1.770 0.340 ;
        RECT  1.770 -0.300 2.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.520 2.820 ;
        RECT  1.520 2.180 1.740 2.820 ;
        RECT  1.740 2.220 2.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.710 0.720 1.870 1.800 ;
        RECT  0.430 0.720 1.710 0.880 ;
        RECT  0.430 1.640 1.710 1.800 ;
        RECT  0.210 1.640 0.430 2.060 ;
    END
END OR4D1

MACRO OR4D2
    CLASS CORE ;
    FOREIGN OR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.960 1.950 2.100 ;
        RECT  1.950 1.390 2.010 2.100 ;
        RECT  1.950 0.420 2.010 0.900 ;
        RECT  2.010 0.420 2.110 2.100 ;
        RECT  2.110 1.960 2.140 2.100 ;
        RECT  2.110 0.780 2.150 1.515 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.005 0.550 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.710 1.005 0.870 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.030 1.005 1.190 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.360 1.005 1.520 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.130 0.300 ;
        RECT  0.130 -0.300 0.350 0.340 ;
        RECT  0.350 -0.300 0.795 0.300 ;
        RECT  0.795 -0.300 1.015 0.340 ;
        RECT  1.015 -0.300 1.510 0.300 ;
        RECT  1.510 -0.300 1.730 0.340 ;
        RECT  1.730 -0.300 2.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.510 2.820 ;
        RECT  1.510 2.180 1.730 2.820 ;
        RECT  1.730 2.220 2.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.830 1.050 1.870 1.270 ;
        RECT  1.710 0.720 1.830 1.800 ;
        RECT  0.430 0.720 1.710 0.880 ;
        RECT  0.430 1.640 1.710 1.800 ;
        RECT  0.210 1.640 0.430 2.060 ;
    END
END OR4D2

MACRO OR4D4
    CLASS CORE ;
    FOREIGN OR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.640 3.470 2.020 ;
        RECT  3.210 0.500 3.470 0.880 ;
        RECT  3.470 0.500 3.890 2.020 ;
        RECT  3.890 1.640 4.250 2.020 ;
        RECT  3.890 0.500 4.250 0.880 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.030 1.090 1.515 ;
        RECT  1.090 1.395 1.990 1.515 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.080 0.670 1.240 ;
        RECT  0.670 1.080 0.790 1.755 ;
        RECT  0.790 1.635 2.310 1.755 ;
        RECT  2.310 1.005 2.470 1.755 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.270 0.765 0.430 1.290 ;
        RECT  0.430 0.765 2.640 0.885 ;
        RECT  2.640 0.765 2.790 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.620 0.300 ;
        RECT  3.620 -0.300 3.840 0.340 ;
        RECT  3.840 -0.300 4.440 0.300 ;
        RECT  4.440 -0.300 4.660 0.340 ;
        RECT  4.660 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.800 2.820 ;
        RECT  2.800 2.180 3.020 2.820 ;
        RECT  3.020 2.220 3.620 2.820 ;
        RECT  3.620 2.180 3.840 2.820 ;
        RECT  3.840 2.220 4.440 2.820 ;
        RECT  4.440 2.180 4.660 2.820 ;
        RECT  4.660 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.030 1.080 3.255 1.240 ;
        RECT  2.910 0.470 3.030 2.050 ;
        RECT  0.400 0.470 2.910 0.630 ;
        RECT  1.410 1.890 2.910 2.050 ;
        LAYER M1 ;
        RECT  3.210 0.500 3.255 0.880 ;
        RECT  3.210 1.640 3.255 2.020 ;
        RECT  4.105 0.500 4.250 0.880 ;
        RECT  4.105 1.640 4.250 2.020 ;
    END
END OR4D4

MACRO OR4D8
    CLASS CORE ;
    FOREIGN OR4D8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  3.150 1.640 4.110 2.020 ;
        RECT  3.180 0.500 4.110 0.880 ;
        RECT  4.110 0.500 4.530 2.020 ;
        RECT  4.530 1.640 5.610 2.020 ;
        RECT  4.530 0.500 5.610 0.880 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.005 1.830 1.235 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.990 1.030 1.150 1.515 ;
        RECT  1.150 1.395 1.990 1.515 ;
        RECT  1.990 1.005 2.150 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.080 0.740 1.240 ;
        RECT  0.740 1.080 0.860 1.755 ;
        RECT  0.860 1.635 2.310 1.755 ;
        RECT  2.310 1.005 2.470 1.755 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.290 0.765 0.450 1.290 ;
        RECT  0.450 0.765 2.640 0.885 ;
        RECT  2.640 0.765 2.790 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.030 1.080 3.770 1.240 ;
        RECT  2.910 0.470 3.030 2.050 ;
        RECT  0.400 0.470 2.910 0.630 ;
        RECT  1.410 1.890 2.910 2.050 ;
        LAYER M1 ;
        RECT  3.150 1.640 3.895 2.020 ;
        RECT  3.180 0.500 3.895 0.880 ;
        RECT  4.745 0.500 5.610 0.880 ;
        RECT  4.745 1.640 5.610 2.020 ;
    END
END OR4D8

MACRO SDF4CQD1
    CLASS CORE ;
    FOREIGN SDF4CQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.350 1.960 8.380 2.100 ;
        RECT  8.380 1.390 8.410 2.100 ;
        RECT  8.380 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.550 2.100 ;
        RECT  8.550 1.960 8.570 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.880 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        RECT  2.470 1.075 2.710 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 3.915 0.300 ;
        RECT  3.915 -0.300 4.135 0.460 ;
        RECT  4.135 -0.300 5.820 0.300 ;
        RECT  5.820 -0.300 6.040 0.740 ;
        RECT  6.040 -0.300 7.300 0.300 ;
        RECT  7.300 -0.300 7.520 0.340 ;
        RECT  7.520 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 5.830 2.820 ;
        RECT  5.830 2.000 6.050 2.820 ;
        RECT  6.050 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.500 0.720 4.640 1.240 ;
        RECT  4.640 1.080 4.855 1.240 ;
        RECT  3.450 1.410 3.580 1.570 ;
        RECT  3.555 0.820 3.580 0.940 ;
        RECT  3.580 0.820 3.700 1.570 ;
        RECT  3.700 1.080 4.190 1.240 ;
        RECT  3.075 0.710 3.185 0.930 ;
        RECT  3.185 0.710 3.305 1.570 ;
        RECT  3.305 1.080 3.320 1.570 ;
        RECT  3.320 1.080 3.455 1.240 ;
        RECT  2.560 1.410 2.835 1.570 ;
        RECT  2.280 0.710 2.835 0.870 ;
        RECT  2.835 0.710 2.955 1.570 ;
        RECT  2.955 1.050 3.045 1.270 ;
        RECT  1.480 0.710 1.770 0.870 ;
        RECT  1.480 1.650 1.860 1.810 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.080 0.880 ;
        RECT  1.080 0.760 1.240 1.420 ;
        RECT  4.470 1.080 4.500 1.240 ;
        RECT  4.820 1.420 4.980 2.050 ;
        RECT  4.820 0.470 4.980 0.820 ;
        RECT  4.375 0.470 4.820 0.590 ;
        RECT  4.255 0.470 4.375 0.700 ;
        RECT  3.795 0.580 4.255 0.700 ;
        RECT  3.675 0.470 3.795 0.700 ;
        RECT  1.350 0.470 3.675 0.590 ;
        RECT  6.030 1.100 6.190 1.510 ;
        RECT  5.360 1.390 6.030 1.510 ;
        RECT  6.390 0.860 6.450 1.790 ;
        RECT  6.330 0.700 6.390 1.790 ;
        RECT  6.230 0.700 6.330 0.980 ;
        RECT  6.210 1.630 6.330 1.790 ;
        RECT  5.850 0.860 6.230 0.980 ;
        RECT  7.010 1.340 7.080 1.750 ;
        RECT  6.920 0.470 7.010 1.750 ;
        RECT  6.890 0.470 6.920 1.460 ;
        RECT  6.670 0.470 6.890 0.590 ;
        RECT  7.600 1.050 7.680 1.270 ;
        RECT  7.480 1.050 7.600 1.510 ;
        RECT  7.450 1.390 7.480 1.510 ;
        RECT  7.330 1.390 7.450 2.050 ;
        RECT  6.800 1.930 7.330 2.050 ;
        RECT  6.770 1.570 6.800 2.050 ;
        RECT  6.640 0.710 6.770 2.050 ;
        RECT  7.920 1.080 8.290 1.240 ;
        RECT  7.880 0.450 7.920 1.510 ;
        RECT  7.880 1.960 7.910 2.100 ;
        RECT  7.800 0.450 7.880 2.100 ;
        RECT  7.700 0.450 7.800 0.870 ;
        RECT  7.720 1.390 7.800 2.100 ;
        RECT  7.690 1.960 7.720 2.100 ;
        RECT  7.340 0.710 7.700 0.870 ;
        RECT  6.610 0.710 6.640 1.690 ;
        RECT  6.450 0.420 6.670 0.590 ;
        RECT  5.690 0.860 5.850 1.270 ;
        RECT  5.200 0.560 5.360 1.670 ;
        RECT  1.110 0.430 1.350 0.590 ;
        RECT  1.200 1.930 4.820 2.050 ;
        RECT  4.310 1.080 4.470 1.620 ;
        RECT  3.425 0.720 3.555 0.940 ;
        RECT  2.700 1.690 4.140 1.810 ;
        RECT  3.080 1.410 3.185 1.570 ;
        RECT  2.340 1.410 2.560 1.810 ;
        RECT  1.360 0.710 1.480 1.810 ;
        RECT  7.180 0.710 7.340 1.270 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDF4CQD1

MACRO SDF4CQD2
    CLASS CORE ;
    FOREIGN SDF4CQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.320 1.960 8.350 2.100 ;
        RECT  8.350 1.390 8.520 2.100 ;
        RECT  8.350 0.420 8.520 0.900 ;
        RECT  8.520 1.960 8.540 2.100 ;
        RECT  8.520 1.390 8.730 1.515 ;
        RECT  8.520 0.780 8.730 0.900 ;
        RECT  8.730 0.780 8.870 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.880 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        RECT  2.470 1.075 2.710 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 3.915 0.300 ;
        RECT  3.915 -0.300 4.135 0.460 ;
        RECT  4.135 -0.300 5.820 0.300 ;
        RECT  5.820 -0.300 6.040 0.740 ;
        RECT  6.040 -0.300 7.220 0.300 ;
        RECT  7.220 -0.300 7.440 0.340 ;
        RECT  7.440 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 5.830 2.820 ;
        RECT  5.830 2.000 6.050 2.820 ;
        RECT  6.050 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.075 0.710 3.185 0.930 ;
        RECT  3.185 0.710 3.305 1.570 ;
        RECT  3.305 1.080 3.320 1.570 ;
        RECT  3.320 1.080 3.455 1.240 ;
        RECT  2.560 1.410 2.835 1.570 ;
        RECT  2.280 0.710 2.835 0.870 ;
        RECT  2.835 0.710 2.955 1.570 ;
        RECT  2.955 1.050 3.045 1.270 ;
        RECT  1.480 0.710 1.770 0.870 ;
        RECT  1.480 1.650 1.860 1.810 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.080 0.880 ;
        RECT  1.080 0.760 1.240 1.420 ;
        RECT  3.900 1.410 4.120 1.810 ;
        RECT  3.700 1.080 4.210 1.240 ;
        RECT  3.580 0.820 3.700 1.570 ;
        RECT  3.555 0.820 3.580 0.940 ;
        RECT  3.450 1.410 3.580 1.570 ;
        RECT  4.640 1.080 4.855 1.240 ;
        RECT  4.500 0.720 4.640 1.240 ;
        RECT  4.380 1.080 4.500 1.810 ;
        RECT  4.820 1.420 4.980 2.050 ;
        RECT  4.820 0.470 4.980 0.820 ;
        RECT  4.375 0.470 4.820 0.590 ;
        RECT  4.255 0.470 4.375 0.700 ;
        RECT  3.795 0.580 4.255 0.700 ;
        RECT  3.675 0.470 3.795 0.700 ;
        RECT  1.350 0.470 3.675 0.590 ;
        RECT  6.030 1.100 6.190 1.510 ;
        RECT  5.360 1.390 6.030 1.510 ;
        RECT  6.390 0.860 6.450 1.790 ;
        RECT  6.330 0.700 6.390 1.790 ;
        RECT  6.230 0.700 6.330 0.980 ;
        RECT  6.210 1.630 6.330 1.790 ;
        RECT  5.850 0.860 6.230 0.980 ;
        RECT  6.890 0.470 7.020 1.750 ;
        RECT  6.670 0.470 6.890 0.590 ;
        RECT  6.860 1.510 6.890 1.750 ;
        RECT  7.540 1.050 7.660 1.270 ;
        RECT  7.420 1.050 7.540 1.510 ;
        RECT  7.330 1.390 7.420 1.510 ;
        RECT  7.210 1.390 7.330 2.050 ;
        RECT  6.830 1.930 7.210 2.050 ;
        RECT  6.730 1.890 6.830 2.050 ;
        RECT  6.730 0.710 6.770 0.930 ;
        RECT  7.900 1.080 8.470 1.240 ;
        RECT  7.830 0.710 7.900 1.510 ;
        RECT  7.780 0.710 7.830 1.890 ;
        RECT  7.300 0.710 7.780 0.870 ;
        RECT  7.660 1.390 7.780 1.890 ;
        RECT  6.610 0.710 6.730 2.050 ;
        RECT  6.450 0.420 6.670 0.590 ;
        RECT  5.690 0.860 5.850 1.270 ;
        RECT  5.200 0.560 5.360 1.670 ;
        RECT  1.110 0.430 1.350 0.590 ;
        RECT  1.200 1.930 4.820 2.050 ;
        RECT  4.280 1.410 4.380 1.810 ;
        RECT  3.425 0.720 3.555 0.940 ;
        RECT  2.700 1.690 3.900 1.810 ;
        RECT  3.080 1.410 3.185 1.570 ;
        RECT  2.340 1.410 2.560 1.810 ;
        RECT  1.360 0.710 1.480 1.810 ;
        RECT  7.140 0.710 7.300 1.230 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDF4CQD2

MACRO SDF4CQD4
    CLASS CORE ;
    FOREIGN SDF4CQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.650 8.590 2.030 ;
        RECT  8.270 0.490 8.590 0.870 ;
        RECT  8.590 0.490 9.010 2.030 ;
        RECT  9.010 1.650 9.180 2.030 ;
        RECT  9.010 0.490 9.180 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 1.830 1.515 ;
        RECT  1.830 1.050 1.880 1.270 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        RECT  2.470 1.080 2.660 1.235 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 3.865 0.300 ;
        RECT  3.865 -0.300 4.085 0.460 ;
        RECT  4.085 -0.300 5.770 0.300 ;
        RECT  5.770 -0.300 5.990 0.740 ;
        RECT  5.990 -0.300 7.170 0.300 ;
        RECT  7.170 -0.300 7.390 0.340 ;
        RECT  7.390 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 5.780 2.820 ;
        RECT  5.780 2.000 6.000 2.820 ;
        RECT  6.000 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.505 0.820 3.530 0.940 ;
        RECT  3.530 0.820 3.650 1.570 ;
        RECT  3.650 1.080 4.160 1.240 ;
        RECT  3.850 1.410 4.070 1.810 ;
        RECT  3.025 0.710 3.135 0.930 ;
        RECT  3.135 0.710 3.255 1.570 ;
        RECT  3.255 1.080 3.270 1.570 ;
        RECT  3.270 1.080 3.405 1.240 ;
        RECT  2.510 1.410 2.785 1.570 ;
        RECT  2.230 0.710 2.785 0.870 ;
        RECT  2.785 0.710 2.905 1.570 ;
        RECT  2.905 1.050 2.995 1.270 ;
        RECT  1.480 0.710 1.770 0.870 ;
        RECT  1.480 1.650 1.860 1.810 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.080 0.880 ;
        RECT  1.080 0.760 1.240 1.420 ;
        RECT  3.400 1.410 3.530 1.570 ;
        RECT  4.590 1.080 4.805 1.240 ;
        RECT  4.450 0.720 4.590 1.240 ;
        RECT  4.330 1.080 4.450 1.810 ;
        RECT  4.770 1.420 4.930 2.050 ;
        RECT  4.770 0.470 4.930 0.820 ;
        RECT  4.325 0.470 4.770 0.590 ;
        RECT  4.205 0.470 4.325 0.700 ;
        RECT  3.745 0.580 4.205 0.700 ;
        RECT  3.625 0.470 3.745 0.700 ;
        RECT  1.350 0.470 3.625 0.590 ;
        RECT  5.980 1.100 6.140 1.510 ;
        RECT  5.310 1.390 5.980 1.510 ;
        RECT  6.340 0.860 6.400 1.790 ;
        RECT  6.280 0.700 6.340 1.790 ;
        RECT  6.180 0.700 6.280 0.980 ;
        RECT  6.160 1.630 6.280 1.790 ;
        RECT  5.800 0.860 6.180 0.980 ;
        RECT  6.840 0.470 6.970 1.750 ;
        RECT  6.620 0.470 6.840 0.590 ;
        RECT  6.810 1.510 6.840 1.750 ;
        RECT  7.490 1.050 7.610 1.270 ;
        RECT  7.370 1.050 7.490 1.510 ;
        RECT  7.280 1.390 7.370 1.510 ;
        RECT  7.160 1.390 7.280 2.050 ;
        RECT  6.780 1.930 7.160 2.050 ;
        RECT  6.680 1.890 6.780 2.050 ;
        RECT  6.680 0.710 6.720 0.930 ;
        RECT  7.850 1.080 8.375 1.240 ;
        RECT  7.790 0.710 7.850 1.510 ;
        RECT  7.770 1.960 7.800 2.100 ;
        RECT  7.770 0.450 7.790 1.510 ;
        RECT  7.730 0.450 7.770 2.100 ;
        RECT  7.570 0.450 7.730 0.870 ;
        RECT  7.610 1.390 7.730 2.100 ;
        RECT  7.580 1.960 7.610 2.100 ;
        RECT  7.250 0.710 7.570 0.870 ;
        RECT  7.090 0.710 7.250 1.230 ;
        RECT  6.560 0.710 6.680 2.050 ;
        RECT  6.400 0.420 6.620 0.590 ;
        RECT  5.640 0.860 5.800 1.270 ;
        RECT  5.150 0.560 5.310 1.670 ;
        RECT  1.110 0.430 1.350 0.590 ;
        RECT  1.200 1.930 4.770 2.050 ;
        RECT  4.230 1.410 4.330 1.810 ;
        RECT  3.375 0.720 3.505 0.940 ;
        RECT  2.650 1.690 3.850 1.810 ;
        RECT  3.030 1.410 3.135 1.570 ;
        RECT  2.290 1.410 2.510 1.810 ;
        RECT  1.360 0.710 1.480 1.810 ;
        RECT  0.100 0.590 0.260 0.880 ;
        LAYER M1 ;
        RECT  8.270 1.650 8.375 2.030 ;
        RECT  8.270 0.490 8.375 0.870 ;
    END
END SDF4CQD4

MACRO SDFCND1
    CLASS CORE ;
    FOREIGN SDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.940 1.940 8.970 2.100 ;
        RECT  8.970 1.390 9.050 2.100 ;
        RECT  8.970 0.420 9.050 0.900 ;
        RECT  9.050 0.420 9.130 2.100 ;
        RECT  9.130 1.940 9.160 2.100 ;
        RECT  9.130 0.760 9.190 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.220 1.960 8.250 2.100 ;
        RECT  8.250 1.390 8.410 2.100 ;
        RECT  8.200 0.710 8.410 0.870 ;
        RECT  8.410 1.960 8.440 2.100 ;
        RECT  8.410 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.285 7.910 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.460 0.300 ;
        RECT  4.460 -0.300 4.610 0.720 ;
        RECT  4.610 -0.300 6.500 0.300 ;
        RECT  6.500 -0.300 6.720 0.590 ;
        RECT  6.720 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.940 2.820 ;
        RECT  4.940 2.040 5.160 2.820 ;
        RECT  5.160 2.220 6.500 2.820 ;
        RECT  6.500 2.180 6.720 2.820 ;
        RECT  6.720 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.810 1.650 7.110 1.810 ;
        RECT  6.810 0.950 7.170 1.070 ;
        RECT  7.170 0.710 7.330 1.070 ;
        RECT  7.330 0.950 7.480 1.070 ;
        RECT  7.480 0.950 7.600 2.050 ;
        RECT  7.600 1.930 7.820 2.050 ;
        RECT  7.600 1.020 8.070 1.160 ;
        RECT  8.070 1.020 8.290 1.180 ;
        RECT  5.510 1.190 5.750 1.310 ;
        RECT  5.750 1.190 5.910 2.050 ;
        RECT  5.910 1.930 7.230 2.050 ;
        RECT  7.190 1.290 7.230 1.530 ;
        RECT  7.230 1.290 7.350 2.050 ;
        RECT  3.850 0.430 3.970 0.960 ;
        RECT  3.970 0.840 4.730 0.960 ;
        RECT  4.730 0.470 4.850 0.960 ;
        RECT  4.850 0.470 5.810 0.610 ;
        RECT  5.810 0.450 6.030 0.610 ;
        RECT  4.310 1.420 5.110 1.580 ;
        RECT  4.970 0.730 5.110 0.950 ;
        RECT  5.110 0.730 5.230 1.580 ;
        RECT  5.230 1.440 5.370 1.580 ;
        RECT  5.370 1.440 5.530 1.960 ;
        RECT  3.610 0.710 3.730 1.910 ;
        RECT  3.730 1.080 3.770 1.910 ;
        RECT  3.770 1.080 4.850 1.200 ;
        RECT  4.850 1.080 4.990 1.300 ;
        RECT  1.410 1.930 3.190 2.050 ;
        RECT  3.190 1.930 3.430 2.090 ;
        RECT  1.340 0.470 3.140 0.590 ;
        RECT  3.140 0.470 3.380 0.630 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  6.670 0.950 6.810 1.810 ;
        RECT  8.850 1.050 8.890 1.290 ;
        RECT  8.710 0.470 8.850 1.290 ;
        RECT  7.000 0.470 8.710 0.590 ;
        RECT  6.880 0.470 7.000 0.830 ;
        RECT  6.330 0.710 6.880 0.830 ;
        RECT  6.170 0.650 6.330 0.975 ;
        RECT  6.170 1.500 6.270 1.720 ;
        RECT  6.160 0.650 6.170 1.720 ;
        RECT  6.030 0.820 6.160 1.720 ;
        RECT  6.310 1.125 6.670 1.345 ;
        RECT  5.350 0.770 5.510 1.310 ;
        RECT  3.700 0.430 3.850 0.590 ;
        RECT  4.090 1.410 4.310 1.580 ;
        RECT  3.570 0.710 3.610 1.195 ;
        RECT  3.940 1.700 4.910 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
        RECT  5.680 0.820 6.030 0.980 ;
    END
END SDFCND1

MACRO SDFCND2
    CLASS CORE ;
    FOREIGN SDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.950 8.990 2.090 ;
        RECT  8.990 1.380 9.150 2.090 ;
        RECT  9.150 1.950 9.180 2.090 ;
        RECT  8.960 0.490 9.180 0.910 ;
        RECT  9.150 1.380 9.370 1.515 ;
        RECT  9.180 0.790 9.370 0.910 ;
        RECT  9.370 0.790 9.510 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.950 8.300 2.090 ;
        RECT  8.300 1.380 8.410 2.090 ;
        RECT  8.240 0.710 8.410 0.870 ;
        RECT  8.410 0.710 8.460 2.090 ;
        RECT  8.460 1.950 8.490 2.090 ;
        RECT  8.460 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.285 7.910 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.460 0.300 ;
        RECT  4.460 -0.300 4.610 0.720 ;
        RECT  4.610 -0.300 6.500 0.300 ;
        RECT  6.500 -0.300 6.720 0.590 ;
        RECT  6.720 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.940 2.820 ;
        RECT  4.940 2.040 5.160 2.820 ;
        RECT  5.160 2.220 6.500 2.820 ;
        RECT  6.500 2.180 6.720 2.820 ;
        RECT  6.720 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.120 1.020 8.290 1.180 ;
        RECT  5.510 1.190 5.750 1.310 ;
        RECT  5.750 1.190 5.910 2.050 ;
        RECT  5.910 1.930 7.230 2.050 ;
        RECT  7.190 1.290 7.230 1.530 ;
        RECT  7.230 1.290 7.350 2.050 ;
        RECT  3.850 0.430 3.970 0.960 ;
        RECT  3.970 0.840 4.730 0.960 ;
        RECT  4.730 0.470 4.850 0.960 ;
        RECT  4.850 0.470 5.810 0.610 ;
        RECT  5.810 0.450 6.050 0.610 ;
        RECT  4.310 1.420 5.110 1.580 ;
        RECT  4.970 0.730 5.110 0.950 ;
        RECT  5.110 0.730 5.230 1.580 ;
        RECT  5.230 1.440 5.370 1.580 ;
        RECT  5.370 1.440 5.530 1.960 ;
        RECT  3.610 0.710 3.730 1.910 ;
        RECT  3.730 1.080 3.770 1.910 ;
        RECT  3.770 1.080 4.850 1.200 ;
        RECT  4.850 1.080 4.990 1.300 ;
        RECT  1.410 1.930 3.190 2.050 ;
        RECT  3.190 1.930 3.430 2.090 ;
        RECT  1.340 0.470 3.140 0.590 ;
        RECT  3.140 0.470 3.380 0.630 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  8.000 0.710 8.120 1.180 ;
        RECT  7.600 0.710 8.000 0.830 ;
        RECT  7.600 1.930 7.820 2.050 ;
        RECT  7.480 0.710 7.600 2.050 ;
        RECT  7.170 0.710 7.480 1.070 ;
        RECT  6.810 0.950 7.170 1.070 ;
        RECT  6.810 1.650 7.110 1.810 ;
        RECT  6.670 0.950 6.810 1.810 ;
        RECT  8.840 1.080 9.080 1.240 ;
        RECT  8.720 0.470 8.840 1.240 ;
        RECT  7.000 0.470 8.720 0.590 ;
        RECT  6.880 0.470 7.000 0.830 ;
        RECT  6.330 0.710 6.880 0.830 ;
        RECT  6.170 0.710 6.330 0.975 ;
        RECT  6.170 1.505 6.270 1.745 ;
        RECT  6.160 0.710 6.170 1.745 ;
        RECT  6.130 0.820 6.160 1.745 ;
        RECT  6.030 0.820 6.130 1.645 ;
        RECT  6.310 1.125 6.670 1.345 ;
        RECT  5.680 0.820 6.030 0.980 ;
        RECT  5.350 0.770 5.510 1.310 ;
        RECT  3.700 0.430 3.850 0.590 ;
        RECT  4.090 1.410 4.310 1.580 ;
        RECT  3.570 0.710 3.610 1.195 ;
        RECT  3.940 1.700 4.910 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
    END
END SDFCND2

MACRO SDFCND4
    CLASS CORE ;
    FOREIGN SDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 1.650 10.830 2.030 ;
        RECT  10.430 0.490 10.830 0.870 ;
        RECT  10.830 0.490 11.250 2.030 ;
        RECT  11.250 1.650 11.360 2.030 ;
        RECT  11.250 0.490 11.360 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.990 1.610 9.230 1.770 ;
        RECT  8.960 0.760 9.230 0.920 ;
        RECT  9.230 0.760 9.650 1.770 ;
        RECT  9.650 1.610 9.960 1.770 ;
        RECT  9.650 0.760 9.960 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 1.190 7.950 1.515 ;
        RECT  7.950 1.285 8.230 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.620 0.720 ;
        RECT  4.620 -0.300 6.510 0.300 ;
        RECT  6.510 -0.300 6.730 0.590 ;
        RECT  6.730 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 8.590 0.300 ;
        RECT  8.590 -0.300 8.810 0.340 ;
        RECT  8.810 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 4.950 2.820 ;
        RECT  4.950 2.040 5.170 2.820 ;
        RECT  5.170 2.220 6.510 2.820 ;
        RECT  6.510 2.180 6.730 2.820 ;
        RECT  6.730 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.200 1.930 3.440 2.090 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  1.410 1.930 3.200 2.050 ;
        RECT  4.860 1.080 5.000 1.300 ;
        RECT  3.780 1.080 4.860 1.200 ;
        RECT  3.740 1.080 3.780 1.910 ;
        RECT  3.620 0.710 3.740 1.910 ;
        RECT  5.380 1.440 5.540 1.960 ;
        RECT  5.240 1.440 5.380 1.580 ;
        RECT  5.120 0.730 5.240 1.580 ;
        RECT  4.980 0.730 5.120 0.950 ;
        RECT  4.320 1.420 5.120 1.580 ;
        RECT  5.820 0.450 6.040 0.610 ;
        RECT  4.860 0.470 5.820 0.610 ;
        RECT  4.740 0.470 4.860 0.960 ;
        RECT  3.980 0.840 4.740 0.960 ;
        RECT  3.860 0.430 3.980 0.960 ;
        RECT  7.250 1.190 7.370 2.050 ;
        RECT  7.210 1.190 7.250 1.410 ;
        RECT  5.920 1.930 7.250 2.050 ;
        RECT  5.760 1.190 5.920 2.050 ;
        RECT  5.520 1.190 5.760 1.310 ;
        RECT  8.560 1.080 8.740 1.240 ;
        RECT  8.440 0.950 8.560 1.240 ;
        RECT  7.610 0.950 8.440 1.070 ;
        RECT  7.610 1.890 7.840 2.050 ;
        RECT  7.490 0.950 7.610 2.050 ;
        RECT  7.340 0.950 7.490 1.070 ;
        RECT  7.180 0.710 7.340 1.070 ;
        RECT  6.820 0.950 7.180 1.070 ;
        RECT  6.820 1.650 7.130 1.810 ;
        RECT  6.680 0.950 6.820 1.810 ;
        RECT  10.260 1.080 10.540 1.240 ;
        RECT  10.140 0.470 10.260 2.050 ;
        RECT  7.010 0.470 10.140 0.590 ;
        RECT  8.220 1.890 10.140 2.050 ;
        RECT  6.890 0.470 7.010 0.830 ;
        RECT  6.340 0.710 6.890 0.830 ;
        RECT  6.180 0.650 6.340 0.975 ;
        RECT  6.180 1.495 6.280 1.715 ;
        RECT  6.170 0.650 6.180 1.715 ;
        RECT  6.040 0.820 6.170 1.715 ;
        RECT  6.320 1.125 6.680 1.345 ;
        RECT  5.360 0.770 5.520 1.310 ;
        RECT  5.690 0.820 6.040 0.980 ;
        RECT  3.710 0.430 3.860 0.590 ;
        RECT  4.100 1.410 4.320 1.580 ;
        RECT  3.580 0.710 3.620 1.195 ;
        RECT  3.950 1.700 4.920 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
        LAYER M1 ;
        RECT  10.430 1.650 10.615 2.030 ;
        RECT  10.430 0.490 10.615 0.870 ;
        RECT  9.865 1.610 9.960 1.770 ;
        RECT  9.865 0.760 9.960 0.920 ;
        RECT  8.990 1.610 9.015 1.770 ;
        RECT  8.960 0.760 9.015 0.920 ;
    END
END SDFCND4

MACRO SDFCNQD1
    CLASS CORE ;
    FOREIGN SDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.720 1.960 7.750 2.100 ;
        RECT  7.750 0.420 7.910 2.100 ;
        RECT  7.910 1.960 7.940 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.130 2.010 1.350 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 6.950 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.620 0.720 ;
        RECT  4.620 -0.300 6.430 0.300 ;
        RECT  6.430 -0.300 6.650 0.490 ;
        RECT  6.650 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.950 2.820 ;
        RECT  4.950 2.040 5.170 2.820 ;
        RECT  5.170 2.220 6.380 2.820 ;
        RECT  6.380 2.180 6.600 2.820 ;
        RECT  6.600 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.230 1.020 7.350 1.470 ;
        RECT  5.920 1.930 7.365 2.050 ;
        RECT  7.350 1.350 7.365 1.470 ;
        RECT  7.365 1.350 7.485 2.050 ;
        RECT  5.930 0.770 6.090 0.980 ;
        RECT  6.090 0.770 6.350 0.930 ;
        RECT  3.860 0.430 3.980 0.960 ;
        RECT  3.980 0.840 4.740 0.960 ;
        RECT  4.740 0.470 4.860 0.960 ;
        RECT  4.860 0.470 5.820 0.610 ;
        RECT  5.820 0.450 6.060 0.610 ;
        RECT  4.320 1.420 5.120 1.580 ;
        RECT  4.980 0.730 5.120 0.950 ;
        RECT  5.120 0.730 5.240 1.580 ;
        RECT  5.240 1.440 5.380 1.580 ;
        RECT  5.380 1.440 5.540 1.960 ;
        RECT  3.620 0.710 3.740 1.910 ;
        RECT  3.740 1.080 3.780 1.910 ;
        RECT  3.780 1.080 4.860 1.200 ;
        RECT  4.860 1.080 5.000 1.300 ;
        RECT  1.410 1.930 3.200 2.050 ;
        RECT  3.200 1.930 3.440 2.090 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.430 ;
        RECT  7.080 1.020 7.230 1.190 ;
        RECT  5.760 1.190 5.920 2.050 ;
        RECT  5.520 1.190 5.760 1.310 ;
        RECT  7.470 0.690 7.630 1.230 ;
        RECT  7.290 0.690 7.470 0.850 ;
        RECT  7.070 0.430 7.290 0.850 ;
        RECT  6.460 1.650 7.190 1.810 ;
        RECT  6.610 0.690 7.070 0.850 ;
        RECT  6.470 0.690 6.610 1.320 ;
        RECT  6.460 1.050 6.470 1.320 ;
        RECT  6.300 1.050 6.460 1.810 ;
        RECT  5.360 0.770 5.520 1.310 ;
        RECT  5.690 0.820 5.930 0.980 ;
        RECT  3.710 0.430 3.860 0.590 ;
        RECT  4.100 1.410 4.320 1.580 ;
        RECT  3.580 0.710 3.620 1.195 ;
        RECT  3.950 1.700 4.920 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
    END
END SDFCNQD1

MACRO SDFCNQD2
    CLASS CORE ;
    FOREIGN SDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.260 1.960 8.290 2.100 ;
        RECT  8.290 1.390 8.410 2.100 ;
        RECT  8.180 0.485 8.410 0.645 ;
        RECT  8.410 0.485 8.450 2.100 ;
        RECT  8.450 1.960 8.480 2.100 ;
        RECT  8.450 0.485 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.130 2.010 1.350 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.190 7.770 1.410 ;
        RECT  7.770 1.005 7.910 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.620 0.720 ;
        RECT  4.620 -0.300 6.430 0.300 ;
        RECT  6.430 -0.300 6.650 0.490 ;
        RECT  6.650 -0.300 7.755 0.300 ;
        RECT  7.755 -0.300 7.975 0.340 ;
        RECT  7.975 -0.300 8.600 0.300 ;
        RECT  8.600 -0.300 8.820 0.340 ;
        RECT  8.820 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.950 2.820 ;
        RECT  4.950 2.040 5.170 2.820 ;
        RECT  5.170 2.220 6.380 2.820 ;
        RECT  6.380 2.180 6.600 2.820 ;
        RECT  6.600 2.220 7.865 2.820 ;
        RECT  7.865 2.180 8.085 2.820 ;
        RECT  8.085 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.430 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.200 1.930 3.440 2.090 ;
        RECT  1.410 1.930 3.200 2.050 ;
        RECT  4.840 1.080 4.980 1.300 ;
        RECT  3.780 1.080 4.840 1.200 ;
        RECT  3.740 1.080 3.780 1.910 ;
        RECT  3.620 0.710 3.740 1.910 ;
        RECT  5.380 1.440 5.540 1.960 ;
        RECT  5.240 1.440 5.380 1.580 ;
        RECT  5.100 0.730 5.240 1.580 ;
        RECT  4.980 0.730 5.100 0.950 ;
        RECT  4.320 1.420 5.100 1.580 ;
        RECT  5.820 0.450 6.060 0.610 ;
        RECT  4.860 0.470 5.820 0.610 ;
        RECT  4.740 0.470 4.860 0.960 ;
        RECT  3.980 0.840 4.740 0.960 ;
        RECT  3.860 0.430 3.980 0.960 ;
        RECT  7.120 1.190 7.240 2.050 ;
        RECT  7.080 1.190 7.120 1.430 ;
        RECT  5.920 1.930 7.120 2.050 ;
        RECT  5.760 1.190 5.920 2.050 ;
        RECT  5.520 1.190 5.760 1.310 ;
        RECT  8.150 1.050 8.280 1.270 ;
        RECT  8.030 0.765 8.150 1.270 ;
        RECT  7.520 0.765 8.030 0.885 ;
        RECT  7.520 1.800 7.710 1.960 ;
        RECT  7.400 0.765 7.520 1.960 ;
        RECT  7.260 0.765 7.400 1.070 ;
        RECT  7.100 0.690 7.260 1.070 ;
        RECT  6.730 0.950 7.100 1.070 ;
        RECT  6.730 1.650 7.000 1.810 ;
        RECT  6.590 0.950 6.730 1.810 ;
        RECT  5.360 0.770 5.520 1.310 ;
        RECT  6.320 1.125 6.590 1.345 ;
        RECT  5.690 0.820 6.370 0.980 ;
        RECT  3.710 0.430 3.860 0.590 ;
        RECT  4.100 1.410 4.320 1.580 ;
        RECT  3.580 0.710 3.620 1.195 ;
        RECT  3.950 1.700 4.920 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
    END
END SDFCNQD2

MACRO SDFCNQD4
    CLASS CORE ;
    FOREIGN SDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.230 1.650 8.590 2.030 ;
        RECT  8.180 0.485 8.590 0.645 ;
        RECT  8.590 0.485 9.010 2.030 ;
        RECT  9.010 1.650 9.160 2.030 ;
        RECT  9.010 0.485 9.180 0.625 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.190 7.770 1.410 ;
        RECT  7.770 1.005 7.910 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.620 0.720 ;
        RECT  4.620 -0.300 6.430 0.300 ;
        RECT  6.430 -0.300 6.650 0.490 ;
        RECT  6.650 -0.300 7.755 0.300 ;
        RECT  7.755 -0.300 7.975 0.340 ;
        RECT  7.975 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 4.950 2.820 ;
        RECT  4.950 2.040 5.170 2.820 ;
        RECT  5.170 2.220 6.380 2.820 ;
        RECT  6.380 2.180 6.600 2.820 ;
        RECT  6.600 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.160 3.260 1.380 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.725 1.630 0.885 ;
        RECT  1.630 0.725 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  3.200 1.930 3.440 2.090 ;
        RECT  1.410 1.930 3.200 2.050 ;
        RECT  4.860 1.080 5.000 1.300 ;
        RECT  3.780 1.080 4.860 1.200 ;
        RECT  3.740 1.080 3.780 1.910 ;
        RECT  3.620 0.710 3.740 1.910 ;
        RECT  5.380 1.440 5.540 1.960 ;
        RECT  5.240 1.440 5.380 1.580 ;
        RECT  5.120 0.730 5.240 1.580 ;
        RECT  4.980 0.730 5.120 0.950 ;
        RECT  4.320 1.420 5.120 1.580 ;
        RECT  5.820 0.450 6.060 0.610 ;
        RECT  4.860 0.470 5.820 0.610 ;
        RECT  4.740 0.470 4.860 0.960 ;
        RECT  3.980 0.840 4.740 0.960 ;
        RECT  3.860 0.430 3.980 0.960 ;
        RECT  7.120 1.190 7.240 2.050 ;
        RECT  7.080 1.190 7.120 1.410 ;
        RECT  5.920 1.930 7.120 2.050 ;
        RECT  5.760 1.190 5.920 2.050 ;
        RECT  5.520 1.190 5.760 1.310 ;
        RECT  8.150 1.080 8.350 1.240 ;
        RECT  8.030 0.765 8.150 1.240 ;
        RECT  7.520 0.765 8.030 0.885 ;
        RECT  7.520 1.800 7.710 1.960 ;
        RECT  7.400 0.765 7.520 1.960 ;
        RECT  7.260 0.765 7.400 1.070 ;
        RECT  7.100 0.690 7.260 1.070 ;
        RECT  6.730 0.950 7.100 1.070 ;
        RECT  6.730 1.650 7.000 1.810 ;
        RECT  6.590 0.950 6.730 1.810 ;
        RECT  6.320 1.125 6.590 1.345 ;
        RECT  5.360 0.770 5.520 1.310 ;
        RECT  5.690 0.820 6.370 0.980 ;
        RECT  3.710 0.430 3.860 0.590 ;
        RECT  4.100 1.410 4.320 1.580 ;
        RECT  3.580 0.710 3.620 1.195 ;
        RECT  3.950 1.700 4.920 1.860 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
        LAYER M1 ;
        RECT  8.230 1.650 8.375 2.030 ;
        RECT  8.180 0.485 8.375 0.645 ;
    END
END SDFCNQD4

MACRO SDFCSND1
    CLASS CORE ;
    FOREIGN SDFCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.725 8.240 1.290 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.600 1.490 8.730 1.650 ;
        RECT  8.630 0.420 8.730 0.910 ;
        RECT  8.730 0.420 8.790 1.650 ;
        RECT  8.790 0.790 8.870 1.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.320 1.960 9.350 2.100 ;
        RECT  9.350 1.390 9.370 2.100 ;
        RECT  9.350 0.420 9.370 0.900 ;
        RECT  9.370 0.420 9.510 2.100 ;
        RECT  9.510 1.960 9.540 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 7.270 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 7.480 0.300 ;
        RECT  7.480 -0.300 7.700 0.340 ;
        RECT  7.700 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.470 2.820 ;
        RECT  2.470 2.180 2.690 2.820 ;
        RECT  2.690 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.760 2.820 ;
        RECT  6.760 1.970 6.980 2.820 ;
        RECT  6.980 2.220 7.560 2.820 ;
        RECT  7.560 2.030 7.780 2.820 ;
        RECT  7.780 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.790 1.080 7.960 1.240 ;
        RECT  7.790 1.770 9.100 1.890 ;
        RECT  9.100 1.030 9.220 1.890 ;
        RECT  9.220 1.030 9.250 1.270 ;
        RECT  6.460 0.470 6.580 1.610 ;
        RECT  6.580 1.450 6.750 1.610 ;
        RECT  6.580 0.470 8.250 0.590 ;
        RECT  7.940 1.490 8.360 1.650 ;
        RECT  8.250 0.430 8.360 0.590 ;
        RECT  8.360 0.430 8.480 1.650 ;
        RECT  8.480 1.050 8.610 1.270 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  6.220 1.160 6.340 2.100 ;
        RECT  6.340 1.730 6.440 2.100 ;
        RECT  6.440 1.730 6.870 1.850 ;
        RECT  6.870 1.490 6.990 1.850 ;
        RECT  6.990 1.490 7.390 1.610 ;
        RECT  7.390 1.030 7.550 1.610 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.940 1.780 6.100 2.090 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.130 3.380 1.350 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.470 1.660 1.710 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  7.670 0.710 7.790 1.890 ;
        RECT  6.790 0.710 7.670 0.870 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  3.690 1.930 3.930 2.100 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.710 ;
        RECT  7.140 1.730 7.670 1.890 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFCSND1

MACRO SDFCSND2
    CLASS CORE ;
    FOREIGN SDFCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.730 1.005 9.190 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.550 1.410 9.690 1.810 ;
        RECT  9.580 0.420 9.690 0.900 ;
        RECT  9.690 0.420 9.740 1.810 ;
        RECT  9.740 0.780 9.770 1.810 ;
        RECT  9.770 0.780 9.830 1.530 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.240 1.940 10.270 2.100 ;
        RECT  10.270 1.390 10.330 2.100 ;
        RECT  10.270 0.420 10.330 0.900 ;
        RECT  10.330 0.420 10.430 2.100 ;
        RECT  10.430 1.940 10.460 2.100 ;
        RECT  10.430 0.780 10.470 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.005 7.910 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 6.970 0.300 ;
        RECT  6.970 -0.300 7.190 0.490 ;
        RECT  7.190 -0.300 9.150 0.300 ;
        RECT  9.150 -0.300 9.370 0.340 ;
        RECT  9.370 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.470 2.820 ;
        RECT  2.470 2.180 2.690 2.820 ;
        RECT  2.690 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.850 2.820 ;
        RECT  6.850 2.030 7.070 2.820 ;
        RECT  7.070 2.220 8.330 2.820 ;
        RECT  8.330 2.010 8.550 2.820 ;
        RECT  8.550 2.220 9.140 2.820 ;
        RECT  9.140 2.180 9.360 2.820 ;
        RECT  9.360 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.940 1.780 6.100 2.100 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.130 3.380 1.350 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.470 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  8.120 1.030 8.280 1.500 ;
        RECT  7.310 1.380 8.120 1.500 ;
        RECT  7.150 1.030 7.310 1.500 ;
        RECT  7.070 1.380 7.150 1.500 ;
        RECT  6.950 1.380 7.070 1.850 ;
        RECT  6.440 1.730 6.950 1.850 ;
        RECT  6.340 1.730 6.440 2.100 ;
        RECT  6.220 1.160 6.340 2.100 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  9.430 1.080 9.570 1.240 ;
        RECT  9.310 0.720 9.430 1.650 ;
        RECT  9.090 0.720 9.310 0.840 ;
        RECT  8.700 1.490 9.310 1.650 ;
        RECT  8.930 0.470 9.090 0.840 ;
        RECT  7.500 0.470 8.930 0.590 ;
        RECT  7.380 0.470 7.500 0.830 ;
        RECT  6.580 0.710 7.380 0.830 ;
        RECT  6.580 1.450 6.750 1.610 ;
        RECT  6.460 0.710 6.580 1.610 ;
        RECT  10.120 1.050 10.210 1.270 ;
        RECT  10.000 1.050 10.120 2.050 ;
        RECT  9.220 1.930 10.000 2.050 ;
        RECT  9.100 1.770 9.220 2.050 ;
        RECT  8.580 1.770 9.100 1.890 ;
        RECT  8.580 1.050 8.610 1.270 ;
        RECT  8.460 0.710 8.580 1.890 ;
        RECT  7.620 0.710 8.460 0.850 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  7.230 1.620 8.460 1.780 ;
        RECT  3.690 1.930 3.930 2.100 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFCSND2

MACRO SDFCSND4
    CLASS CORE ;
    FOREIGN SDFCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.730 0.725 8.870 1.235 ;
        RECT  8.870 1.075 9.005 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.430 1.600 9.870 1.760 ;
        RECT  9.450 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 1.760 ;
        RECT  10.290 0.490 10.360 0.870 ;
        RECT  10.290 1.600 10.380 1.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.830 1.650 11.150 2.030 ;
        RECT  10.830 0.490 11.150 0.870 ;
        RECT  11.150 0.490 11.570 2.030 ;
        RECT  11.570 1.650 11.740 2.030 ;
        RECT  11.570 0.490 11.740 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.005 7.910 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 6.880 0.300 ;
        RECT  6.880 -0.300 7.100 0.490 ;
        RECT  7.100 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.760 2.820 ;
        RECT  6.760 2.030 6.980 2.820 ;
        RECT  6.980 2.220 8.240 2.820 ;
        RECT  8.240 2.010 8.460 2.820 ;
        RECT  8.460 2.220 9.040 2.820 ;
        RECT  9.040 2.180 9.260 2.820 ;
        RECT  9.260 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.130 3.380 1.350 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.470 1.660 1.710 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  5.940 1.780 6.100 2.100 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  8.030 1.030 8.190 1.500 ;
        RECT  7.220 1.380 8.030 1.500 ;
        RECT  7.060 1.030 7.220 1.500 ;
        RECT  6.980 1.380 7.060 1.500 ;
        RECT  6.860 1.380 6.980 1.850 ;
        RECT  6.440 1.730 6.860 1.850 ;
        RECT  6.340 1.730 6.440 2.100 ;
        RECT  6.220 1.160 6.340 2.100 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  9.245 1.080 9.570 1.240 ;
        RECT  9.125 0.430 9.245 1.650 ;
        RECT  8.810 0.430 9.125 0.590 ;
        RECT  8.610 1.490 9.125 1.650 ;
        RECT  7.410 0.470 8.810 0.590 ;
        RECT  7.290 0.470 7.410 0.830 ;
        RECT  6.580 0.710 7.290 0.830 ;
        RECT  6.580 1.450 6.740 1.610 ;
        RECT  6.460 0.710 6.580 1.610 ;
        RECT  10.660 1.050 10.890 1.270 ;
        RECT  10.540 1.050 10.660 2.050 ;
        RECT  9.130 1.930 10.540 2.050 ;
        RECT  9.010 1.770 9.130 2.050 ;
        RECT  8.490 1.770 9.010 1.890 ;
        RECT  8.490 1.050 8.520 1.270 ;
        RECT  8.370 0.710 8.490 1.890 ;
        RECT  7.530 0.710 8.370 0.870 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  7.140 1.620 8.370 1.780 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  3.690 1.930 3.930 2.100 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.710 ;
        RECT  0.080 0.760 0.100 1.850 ;
        LAYER M1 ;
        RECT  10.830 1.650 10.935 2.030 ;
        RECT  10.830 0.490 10.935 0.870 ;
        RECT  9.450 0.490 9.655 0.870 ;
        RECT  9.430 1.600 9.655 1.760 ;
    END
END SDFCSND4

MACRO SDFD1
    CLASS CORE ;
    FOREIGN SDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.720 1.960 7.750 2.100 ;
        RECT  7.750 0.420 7.910 2.100 ;
        RECT  7.910 1.960 7.940 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.890 1.960 6.920 2.100 ;
        RECT  6.920 1.390 7.080 2.100 ;
        RECT  7.080 1.960 7.110 2.100 ;
        RECT  7.080 1.390 7.130 1.515 ;
        RECT  6.920 0.710 7.130 0.870 ;
        RECT  7.130 0.710 7.270 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 2.700 0.300 ;
        RECT  2.700 -0.300 2.920 0.340 ;
        RECT  2.920 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.740 ;
        RECT  4.690 -0.300 6.150 0.300 ;
        RECT  6.150 -0.300 6.370 0.340 ;
        RECT  6.370 -0.300 7.320 0.300 ;
        RECT  7.320 -0.300 7.540 0.340 ;
        RECT  7.540 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.700 2.820 ;
        RECT  2.700 2.180 2.920 2.820 ;
        RECT  2.920 2.220 4.380 2.820 ;
        RECT  4.380 2.000 4.600 2.820 ;
        RECT  4.600 2.220 6.140 2.820 ;
        RECT  6.140 2.180 6.360 2.820 ;
        RECT  6.360 2.220 7.310 2.820 ;
        RECT  7.310 2.180 7.530 2.820 ;
        RECT  7.530 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.800 1.080 7.010 1.240 ;
        RECT  5.260 0.710 5.350 2.050 ;
        RECT  5.350 0.710 5.420 0.930 ;
        RECT  5.350 1.930 6.190 2.050 ;
        RECT  6.190 1.390 6.310 2.050 ;
        RECT  6.310 1.390 6.340 1.510 ;
        RECT  6.340 1.050 6.460 1.510 ;
        RECT  6.460 1.050 6.560 1.270 ;
        RECT  5.470 1.150 5.540 1.750 ;
        RECT  5.320 0.470 5.540 0.590 ;
        RECT  5.540 0.470 5.630 1.750 ;
        RECT  5.630 0.470 5.660 1.270 ;
        RECT  4.500 0.860 4.880 0.980 ;
        RECT  4.760 1.630 4.940 1.790 ;
        RECT  4.880 0.700 4.940 0.980 ;
        RECT  4.940 0.700 5.040 1.790 ;
        RECT  5.040 0.860 5.060 1.790 ;
        RECT  4.010 1.390 4.660 1.510 ;
        RECT  4.660 1.100 4.820 1.510 ;
        RECT  1.350 0.470 3.440 0.590 ;
        RECT  3.440 0.470 3.680 0.630 ;
        RECT  1.410 1.930 3.470 2.050 ;
        RECT  3.470 1.420 3.630 2.050 ;
        RECT  3.150 0.710 3.170 0.930 ;
        RECT  3.170 0.710 3.290 1.810 ;
        RECT  3.290 1.080 3.565 1.240 ;
        RECT  2.280 0.710 2.910 0.870 ;
        RECT  2.910 0.710 3.030 1.810 ;
        RECT  3.030 1.050 3.050 1.270 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.460 1.860 1.620 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  6.740 0.710 6.800 1.510 ;
        RECT  6.740 1.960 6.770 2.100 ;
        RECT  6.680 0.710 6.740 2.100 ;
        RECT  6.200 0.710 6.680 0.870 ;
        RECT  6.580 1.390 6.680 2.100 ;
        RECT  6.550 1.960 6.580 2.100 ;
        RECT  7.470 0.470 7.630 1.290 ;
        RECT  5.920 0.470 7.470 0.590 ;
        RECT  5.910 0.470 5.920 1.580 ;
        RECT  5.780 0.470 5.910 1.810 ;
        RECT  5.750 1.460 5.780 1.810 ;
        RECT  6.040 0.710 6.200 1.270 ;
        RECT  5.190 0.810 5.260 2.050 ;
        RECT  5.100 0.420 5.320 0.590 ;
        RECT  4.340 0.860 4.500 1.270 ;
        RECT  3.850 0.450 4.010 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.150 1.590 3.170 1.810 ;
        RECT  2.350 1.650 2.910 1.810 ;
        RECT  1.530 0.710 1.650 1.620 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFD1

MACRO SDFD2
    CLASS CORE ;
    FOREIGN SDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.000 1.960 8.030 2.100 ;
        RECT  8.030 1.390 8.090 2.100 ;
        RECT  8.030 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.190 2.100 ;
        RECT  8.190 1.960 8.220 2.100 ;
        RECT  8.190 0.780 8.230 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.220 1.960 7.250 2.100 ;
        RECT  7.250 1.390 7.410 2.100 ;
        RECT  7.410 1.960 7.440 2.100 ;
        RECT  7.410 1.390 7.450 1.515 ;
        RECT  7.230 0.710 7.450 0.870 ;
        RECT  7.450 0.710 7.590 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 2.680 0.300 ;
        RECT  2.680 -0.300 2.900 0.340 ;
        RECT  2.900 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.740 ;
        RECT  4.670 -0.300 6.130 0.300 ;
        RECT  6.130 -0.300 6.350 0.340 ;
        RECT  6.350 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.680 2.820 ;
        RECT  2.680 2.180 2.900 2.820 ;
        RECT  2.900 2.220 4.360 2.820 ;
        RECT  4.360 2.000 4.580 2.820 ;
        RECT  4.580 2.220 6.120 2.820 ;
        RECT  6.120 2.180 6.340 2.820 ;
        RECT  6.340 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.420 0.470 3.660 0.630 ;
        RECT  1.410 1.930 3.450 2.050 ;
        RECT  3.450 1.420 3.610 2.050 ;
        RECT  3.130 0.710 3.150 0.930 ;
        RECT  3.150 0.710 3.270 1.810 ;
        RECT  3.270 1.080 3.545 1.240 ;
        RECT  2.280 0.710 2.890 0.870 ;
        RECT  2.890 0.710 3.010 1.810 ;
        RECT  3.010 1.050 3.030 1.270 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.430 1.810 1.670 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  1.350 0.470 3.420 0.590 ;
        RECT  4.640 1.100 4.800 1.510 ;
        RECT  3.990 1.390 4.640 1.510 ;
        RECT  5.020 0.860 5.040 1.790 ;
        RECT  4.920 0.700 5.020 1.790 ;
        RECT  4.860 0.700 4.920 0.980 ;
        RECT  4.740 1.630 4.920 1.790 ;
        RECT  4.480 0.860 4.860 0.980 ;
        RECT  5.610 0.470 5.640 1.270 ;
        RECT  5.520 0.470 5.610 1.750 ;
        RECT  5.300 0.470 5.520 0.590 ;
        RECT  5.450 1.150 5.520 1.750 ;
        RECT  6.440 1.050 6.540 1.270 ;
        RECT  6.320 1.050 6.440 1.510 ;
        RECT  6.290 1.390 6.320 1.510 ;
        RECT  6.170 1.390 6.290 2.050 ;
        RECT  5.330 1.930 6.170 2.050 ;
        RECT  5.330 0.710 5.400 0.930 ;
        RECT  5.240 0.710 5.330 2.050 ;
        RECT  6.780 1.080 7.320 1.240 ;
        RECT  6.720 0.710 6.780 1.700 ;
        RECT  6.660 0.710 6.720 2.080 ;
        RECT  6.180 0.710 6.660 0.870 ;
        RECT  6.560 1.580 6.660 2.080 ;
        RECT  7.750 0.470 7.910 1.290 ;
        RECT  5.900 0.470 7.750 0.590 ;
        RECT  5.890 0.470 5.900 1.580 ;
        RECT  5.760 0.470 5.890 1.810 ;
        RECT  6.020 0.710 6.180 1.270 ;
        RECT  5.730 1.460 5.760 1.810 ;
        RECT  5.170 0.810 5.240 2.050 ;
        RECT  5.080 0.420 5.300 0.590 ;
        RECT  4.320 0.860 4.480 1.270 ;
        RECT  3.830 0.450 3.990 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.130 1.590 3.150 1.810 ;
        RECT  2.350 1.650 2.890 1.810 ;
        RECT  1.530 0.710 1.650 1.575 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFD2

MACRO SDFD4
    CLASS CORE ;
    FOREIGN SDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.560 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.230 1.650 9.550 2.030 ;
        RECT  9.230 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 2.030 ;
        RECT  9.970 1.650 10.140 2.030 ;
        RECT  9.970 0.490 10.140 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.850 1.650 8.270 2.030 ;
        RECT  7.830 0.710 8.270 0.870 ;
        RECT  8.270 0.710 8.690 2.030 ;
        RECT  8.690 1.650 8.760 2.030 ;
        RECT  8.690 0.710 8.780 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.610 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 4.340 0.300 ;
        RECT  4.340 -0.300 4.560 0.740 ;
        RECT  4.560 -0.300 5.960 0.300 ;
        RECT  5.960 -0.300 6.180 0.340 ;
        RECT  6.180 -0.300 6.760 0.300 ;
        RECT  6.760 -0.300 6.980 0.340 ;
        RECT  6.980 -0.300 10.560 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 4.350 2.820 ;
        RECT  4.350 2.030 4.570 2.820 ;
        RECT  4.570 2.220 6.070 2.820 ;
        RECT  6.070 2.180 6.290 2.820 ;
        RECT  6.290 2.220 10.560 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  1.650 1.430 1.810 1.670 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  2.900 1.050 2.920 1.270 ;
        RECT  2.780 0.710 2.900 1.810 ;
        RECT  2.170 0.710 2.780 0.870 ;
        RECT  3.160 1.080 3.435 1.240 ;
        RECT  3.040 0.710 3.160 1.810 ;
        RECT  3.020 0.710 3.040 0.930 ;
        RECT  3.340 1.420 3.500 2.050 ;
        RECT  1.410 1.930 3.340 2.050 ;
        RECT  3.310 0.470 3.550 0.630 ;
        RECT  1.350 0.470 3.310 0.590 ;
        RECT  4.530 1.100 4.690 1.510 ;
        RECT  3.880 1.390 4.530 1.510 ;
        RECT  4.910 0.860 4.970 1.790 ;
        RECT  4.850 0.700 4.910 1.790 ;
        RECT  4.750 0.700 4.850 0.980 ;
        RECT  4.730 1.630 4.850 1.790 ;
        RECT  4.370 0.860 4.750 0.980 ;
        RECT  5.530 1.150 5.600 1.750 ;
        RECT  5.440 0.470 5.530 1.750 ;
        RECT  5.410 0.470 5.440 1.275 ;
        RECT  5.190 0.470 5.410 0.590 ;
        RECT  7.160 1.030 7.320 1.510 ;
        RECT  6.890 1.390 7.160 1.510 ;
        RECT  6.770 1.390 6.890 2.050 ;
        RECT  5.320 1.930 6.770 2.050 ;
        RECT  5.290 1.395 5.320 2.050 ;
        RECT  5.160 0.710 5.290 2.050 ;
        RECT  7.660 1.080 7.955 1.240 ;
        RECT  7.540 0.710 7.660 1.775 ;
        RECT  6.940 0.710 7.540 0.870 ;
        RECT  7.380 1.650 7.540 1.775 ;
        RECT  7.160 1.650 7.380 2.070 ;
        RECT  6.820 0.710 6.940 1.240 ;
        RECT  9.090 1.050 9.270 1.270 ;
        RECT  8.930 0.470 9.090 1.270 ;
        RECT  6.580 0.470 8.930 0.590 ;
        RECT  6.500 1.590 6.640 1.810 ;
        RECT  6.360 0.470 6.580 0.680 ;
        RECT  5.880 1.590 6.500 1.710 ;
        RECT  5.840 0.560 6.360 0.680 ;
        RECT  5.840 1.590 5.880 1.810 ;
        RECT  5.720 0.560 5.840 1.810 ;
        RECT  5.650 0.560 5.720 1.000 ;
        RECT  6.600 1.080 6.820 1.240 ;
        RECT  5.130 0.710 5.160 1.515 ;
        RECT  4.970 0.420 5.190 0.590 ;
        RECT  4.210 0.860 4.370 1.270 ;
        RECT  3.720 0.450 3.880 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.020 1.590 3.040 1.810 ;
        RECT  2.240 1.650 2.780 1.810 ;
        RECT  1.530 0.710 1.650 1.575 ;
        RECT  0.100 0.590 0.260 0.880 ;
        LAYER M1 ;
        RECT  9.230 1.650 9.335 2.030 ;
        RECT  9.230 0.490 9.335 0.870 ;
        RECT  7.850 1.650 8.055 2.030 ;
        RECT  7.830 0.710 8.055 0.870 ;
    END
END SDFD4

MACRO SDFKCND1
    CLASS CORE ;
    FOREIGN SDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.060 1.530 8.090 2.030 ;
        RECT  8.060 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.220 2.030 ;
        RECT  8.220 0.780 8.230 1.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.340 1.530 7.450 1.750 ;
        RECT  7.360 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.520 1.750 ;
        RECT  7.520 0.780 7.590 1.750 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.760 0.300 ;
        RECT  1.760 -0.300 1.980 0.490 ;
        RECT  1.980 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.350 ;
        RECT  3.630 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.830 2.820 ;
        RECT  1.830 2.030 2.050 2.820 ;
        RECT  2.050 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 3.455 2.820 ;
        RECT  3.455 2.160 3.675 2.820 ;
        RECT  3.675 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 6.595 2.820 ;
        RECT  6.595 2.160 6.815 2.820 ;
        RECT  6.815 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.160 0.460 6.280 1.420 ;
        RECT  5.905 1.880 6.435 2.040 ;
        RECT  6.280 1.300 6.435 1.420 ;
        RECT  6.435 1.300 6.555 2.040 ;
        RECT  6.555 1.300 6.775 1.420 ;
        RECT  6.775 1.160 6.935 1.420 ;
        RECT  6.040 1.540 6.140 1.680 ;
        RECT  6.140 1.540 6.295 1.760 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.750 0.540 5.800 0.780 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  4.210 0.450 4.450 0.620 ;
        RECT  3.120 0.720 3.550 0.880 ;
        RECT  3.550 0.720 3.670 1.760 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.590 0.970 2.730 1.490 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  7.875 1.050 7.970 1.270 ;
        RECT  7.755 1.050 7.875 2.050 ;
        RECT  7.200 1.930 7.755 2.050 ;
        RECT  7.080 0.450 7.200 2.050 ;
        RECT  6.960 0.450 7.080 0.610 ;
        RECT  6.615 0.910 7.080 1.030 ;
        RECT  6.925 1.580 7.080 1.740 ;
        RECT  6.455 0.910 6.615 1.180 ;
        RECT  5.970 0.460 6.160 0.620 ;
        RECT  5.880 0.870 6.040 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.090 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
    END
END SDFKCND1

MACRO SDFKCND2
    CLASS CORE ;
    FOREIGN SDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.350 1.530 8.410 2.030 ;
        RECT  8.350 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.510 2.030 ;
        RECT  8.510 0.780 8.550 1.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.590 1.560 7.770 1.720 ;
        RECT  7.660 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.820 1.720 ;
        RECT  7.820 0.780 7.910 1.720 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.760 0.300 ;
        RECT  1.760 -0.300 1.980 0.490 ;
        RECT  1.980 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.350 ;
        RECT  3.630 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.830 2.820 ;
        RECT  1.830 2.030 2.050 2.820 ;
        RECT  2.050 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 3.455 2.820 ;
        RECT  3.455 2.160 3.675 2.820 ;
        RECT  3.675 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 6.595 2.820 ;
        RECT  6.595 2.160 6.815 2.820 ;
        RECT  6.815 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  4.210 0.450 4.450 0.620 ;
        RECT  3.120 0.720 3.550 0.880 ;
        RECT  3.550 0.720 3.670 1.760 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.590 0.970 2.730 1.490 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  5.750 0.540 5.800 0.780 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  6.140 1.540 6.295 1.760 ;
        RECT  6.040 1.540 6.140 1.680 ;
        RECT  6.775 1.160 6.935 1.420 ;
        RECT  6.555 1.300 6.775 1.420 ;
        RECT  6.435 1.300 6.555 2.040 ;
        RECT  6.280 1.300 6.435 1.420 ;
        RECT  5.905 1.880 6.435 2.040 ;
        RECT  6.160 0.460 6.280 1.420 ;
        RECT  8.175 1.050 8.270 1.270 ;
        RECT  8.055 1.050 8.175 2.050 ;
        RECT  7.200 1.930 8.055 2.050 ;
        RECT  7.080 0.450 7.200 2.050 ;
        RECT  6.960 0.450 7.080 0.610 ;
        RECT  6.615 0.910 7.080 1.030 ;
        RECT  6.925 1.580 7.080 1.740 ;
        RECT  6.455 0.910 6.615 1.180 ;
        RECT  5.970 0.460 6.160 0.620 ;
        RECT  5.880 0.870 6.040 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.090 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
    END
END SDFKCND2

MACRO SDFKCND4
    CLASS CORE ;
    FOREIGN SDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.170 1.650 10.510 2.030 ;
        RECT  10.190 0.490 10.510 0.870 ;
        RECT  10.510 0.490 10.930 2.030 ;
        RECT  10.930 1.650 11.100 2.030 ;
        RECT  10.930 0.490 11.100 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.770 1.560 8.910 1.720 ;
        RECT  8.810 0.490 8.910 0.870 ;
        RECT  8.910 0.490 9.330 1.720 ;
        RECT  9.330 1.560 9.720 1.720 ;
        RECT  9.330 0.490 9.720 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.760 0.300 ;
        RECT  1.760 -0.300 1.980 0.490 ;
        RECT  1.980 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 6.010 0.300 ;
        RECT  6.010 -0.300 6.230 0.740 ;
        RECT  6.230 -0.300 11.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.780 2.820 ;
        RECT  1.780 2.030 2.000 2.820 ;
        RECT  2.000 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 5.925 2.820 ;
        RECT  5.925 1.760 6.145 2.820 ;
        RECT  6.145 2.220 7.775 2.820 ;
        RECT  7.775 2.160 7.995 2.820 ;
        RECT  7.995 2.220 11.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.590 0.970 2.730 1.490 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  3.550 0.720 3.670 1.760 ;
        RECT  3.120 0.720 3.550 0.880 ;
        RECT  4.210 0.470 4.450 0.630 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  6.915 0.720 6.940 0.940 ;
        RECT  6.800 0.720 6.915 1.760 ;
        RECT  6.755 0.860 6.800 1.760 ;
        RECT  5.800 0.860 6.755 0.980 ;
        RECT  5.750 0.540 5.800 0.980 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  7.320 1.540 7.475 1.760 ;
        RECT  7.230 1.540 7.320 1.680 ;
        RECT  7.955 1.160 8.115 1.420 ;
        RECT  7.735 1.300 7.955 1.420 ;
        RECT  7.615 1.300 7.735 2.040 ;
        RECT  7.470 1.300 7.615 1.420 ;
        RECT  6.535 1.880 7.615 2.040 ;
        RECT  7.350 0.470 7.470 1.420 ;
        RECT  7.170 0.470 7.350 0.620 ;
        RECT  6.590 0.470 7.170 0.600 ;
        RECT  6.350 0.470 6.590 0.630 ;
        RECT  10.045 1.050 10.230 1.270 ;
        RECT  9.925 1.050 10.045 2.050 ;
        RECT  8.380 1.930 9.925 2.050 ;
        RECT  8.260 0.450 8.380 2.050 ;
        RECT  8.140 0.450 8.260 0.610 ;
        RECT  7.795 0.910 8.260 1.030 ;
        RECT  8.105 1.580 8.260 1.740 ;
        RECT  7.635 0.910 7.795 1.180 ;
        RECT  6.375 1.540 6.535 2.040 ;
        RECT  7.070 0.870 7.230 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.090 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
        LAYER M1 ;
        RECT  10.190 0.490 10.295 0.870 ;
        RECT  10.170 1.650 10.295 2.030 ;
        RECT  9.545 1.560 9.720 1.720 ;
        RECT  9.545 0.490 9.720 0.870 ;
    END
END SDFKCND4

MACRO SDFKCNQD1
    CLASS CORE ;
    FOREIGN SDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.310 1.950 7.340 2.090 ;
        RECT  7.340 1.380 7.450 2.090 ;
        RECT  7.390 0.420 7.450 0.900 ;
        RECT  7.450 0.420 7.500 2.090 ;
        RECT  7.500 1.950 7.530 2.090 ;
        RECT  7.500 0.420 7.550 1.515 ;
        RECT  7.550 0.780 7.590 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.710 0.300 ;
        RECT  1.710 -0.300 1.930 0.490 ;
        RECT  1.930 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.350 ;
        RECT  3.630 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.780 2.820 ;
        RECT  1.780 2.030 2.000 2.820 ;
        RECT  2.000 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 3.455 2.820 ;
        RECT  3.455 2.160 3.675 2.820 ;
        RECT  3.675 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 6.595 2.820 ;
        RECT  6.595 2.160 6.815 2.820 ;
        RECT  6.815 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  4.210 0.470 4.450 0.630 ;
        RECT  3.120 0.725 3.550 0.885 ;
        RECT  3.550 0.725 3.670 1.760 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.590 0.980 2.730 1.490 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  5.750 0.540 5.800 0.780 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  6.140 1.540 6.295 1.760 ;
        RECT  6.040 1.540 6.140 1.680 ;
        RECT  6.765 1.160 6.945 1.420 ;
        RECT  6.555 1.300 6.765 1.420 ;
        RECT  6.435 1.300 6.555 2.040 ;
        RECT  6.280 1.300 6.435 1.420 ;
        RECT  5.905 1.880 6.435 2.040 ;
        RECT  6.160 0.460 6.280 1.420 ;
        RECT  7.070 0.420 7.190 1.740 ;
        RECT  7.030 0.420 7.070 1.030 ;
        RECT  6.925 1.580 7.070 1.740 ;
        RECT  6.615 0.910 7.030 1.030 ;
        RECT  5.970 0.460 6.160 0.620 ;
        RECT  5.880 0.870 6.040 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.100 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
        RECT  6.455 0.910 6.615 1.180 ;
    END
END SDFKCNQD1

MACRO SDFKCNQD2
    CLASS CORE ;
    FOREIGN SDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.610 1.950 7.640 2.090 ;
        RECT  7.640 1.380 7.770 2.090 ;
        RECT  7.660 0.420 7.770 0.900 ;
        RECT  7.770 0.420 7.800 2.090 ;
        RECT  7.800 0.420 7.820 1.515 ;
        RECT  7.800 1.950 7.830 2.090 ;
        RECT  7.820 0.780 7.910 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.710 0.300 ;
        RECT  1.710 -0.300 1.930 0.490 ;
        RECT  1.930 -0.300 3.410 0.300 ;
        RECT  3.410 -0.300 3.630 0.350 ;
        RECT  3.630 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.780 2.820 ;
        RECT  1.780 2.030 2.000 2.820 ;
        RECT  2.000 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 3.455 2.820 ;
        RECT  3.455 2.160 3.675 2.820 ;
        RECT  3.675 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 6.595 2.820 ;
        RECT  6.595 2.160 6.815 2.820 ;
        RECT  6.815 2.220 7.210 2.820 ;
        RECT  7.210 2.180 7.430 2.820 ;
        RECT  7.430 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  4.210 0.470 4.450 0.630 ;
        RECT  3.120 0.720 3.550 0.880 ;
        RECT  3.550 0.720 3.670 1.760 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.590 0.970 2.730 1.490 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  5.750 0.540 5.800 0.780 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  6.140 1.540 6.295 1.760 ;
        RECT  6.040 1.540 6.140 1.680 ;
        RECT  6.775 1.160 6.935 1.420 ;
        RECT  6.555 1.300 6.775 1.420 ;
        RECT  6.435 1.300 6.555 2.040 ;
        RECT  6.280 1.300 6.435 1.420 ;
        RECT  5.905 1.880 6.435 2.040 ;
        RECT  6.160 0.460 6.280 1.420 ;
        RECT  7.080 0.450 7.200 1.740 ;
        RECT  6.960 0.450 7.080 0.610 ;
        RECT  6.615 0.910 7.080 1.030 ;
        RECT  6.925 1.580 7.080 1.740 ;
        RECT  5.970 0.460 6.160 0.620 ;
        RECT  5.880 0.870 6.040 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.100 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
        RECT  6.455 0.910 6.615 1.180 ;
    END
END SDFKCNQD2

MACRO SDFKCNQD4
    CLASS CORE ;
    FOREIGN SDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.850 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.210 1.000 2.330 1.220 ;
        RECT  2.330 0.725 2.470 1.235 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.790 1.650 9.230 2.030 ;
        RECT  8.810 0.490 9.230 0.870 ;
        RECT  9.230 0.490 9.650 2.030 ;
        RECT  9.650 1.650 9.700 2.030 ;
        RECT  9.650 0.490 9.720 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.005 3.430 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.410 0.725 0.550 1.300 ;
        RECT  0.550 1.140 0.770 1.300 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.710 0.300 ;
        RECT  1.710 -0.300 1.930 0.490 ;
        RECT  1.930 -0.300 5.230 0.300 ;
        RECT  5.230 -0.300 5.450 0.760 ;
        RECT  5.450 -0.300 6.010 0.300 ;
        RECT  6.010 -0.300 6.230 0.740 ;
        RECT  6.230 -0.300 9.890 0.300 ;
        RECT  9.890 -0.300 10.110 0.340 ;
        RECT  10.110 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.780 2.820 ;
        RECT  1.780 2.030 2.000 2.820 ;
        RECT  2.000 2.220 2.385 2.820 ;
        RECT  2.385 2.160 2.605 2.820 ;
        RECT  2.605 2.220 5.165 2.820 ;
        RECT  5.165 1.760 5.385 2.820 ;
        RECT  5.385 2.220 5.925 2.820 ;
        RECT  5.925 1.760 6.145 2.820 ;
        RECT  6.145 2.220 7.775 2.820 ;
        RECT  7.775 2.160 7.995 2.820 ;
        RECT  7.995 2.220 8.390 2.820 ;
        RECT  8.390 2.160 8.610 2.820 ;
        RECT  8.610 2.220 9.880 2.820 ;
        RECT  9.880 2.180 10.100 2.820 ;
        RECT  10.100 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.250 1.930 0.780 2.050 ;
        RECT  0.710 0.420 0.870 1.010 ;
        RECT  0.780 1.570 0.890 2.050 ;
        RECT  0.870 0.890 0.890 1.010 ;
        RECT  0.890 0.890 0.940 2.050 ;
        RECT  0.940 0.890 1.010 1.690 ;
        RECT  2.090 1.360 2.320 1.520 ;
        RECT  2.090 0.660 2.210 0.880 ;
        RECT  1.970 0.660 2.090 1.520 ;
        RECT  1.530 1.365 1.970 1.520 ;
        RECT  2.590 0.970 2.730 1.490 ;
        RECT  2.575 1.370 2.590 1.490 ;
        RECT  2.455 1.370 2.575 1.890 ;
        RECT  1.250 1.730 2.455 1.890 ;
        RECT  1.130 0.530 1.250 1.890 ;
        RECT  3.670 1.050 3.835 1.270 ;
        RECT  3.550 0.720 3.670 1.760 ;
        RECT  3.120 0.720 3.550 0.880 ;
        RECT  4.210 0.470 4.450 0.630 ;
        RECT  4.135 1.890 4.375 2.050 ;
        RECT  2.985 0.470 4.210 0.590 ;
        RECT  3.005 1.890 4.135 2.010 ;
        RECT  2.985 1.640 3.005 2.070 ;
        RECT  2.940 0.470 2.985 2.070 ;
        RECT  2.860 0.430 2.940 2.070 ;
        RECT  2.720 0.430 2.860 0.850 ;
        RECT  4.105 1.130 4.505 1.290 ;
        RECT  3.985 0.740 4.105 1.660 ;
        RECT  3.790 0.740 3.985 0.900 ;
        RECT  5.340 0.900 5.500 1.300 ;
        RECT  4.780 0.900 5.340 1.020 ;
        RECT  4.755 0.590 4.780 1.020 ;
        RECT  4.635 0.590 4.755 1.920 ;
        RECT  4.620 0.590 4.635 0.830 ;
        RECT  6.915 0.720 6.940 0.940 ;
        RECT  6.800 0.720 6.915 1.760 ;
        RECT  6.755 0.860 6.800 1.760 ;
        RECT  5.800 0.860 6.755 0.980 ;
        RECT  5.750 0.540 5.800 0.980 ;
        RECT  5.630 0.540 5.750 1.980 ;
        RECT  5.575 1.460 5.630 1.980 ;
        RECT  5.190 1.460 5.575 1.580 ;
        RECT  5.060 1.150 5.190 1.580 ;
        RECT  7.320 1.540 7.475 1.760 ;
        RECT  7.230 1.540 7.320 1.680 ;
        RECT  7.955 1.160 8.115 1.420 ;
        RECT  7.735 1.300 7.955 1.420 ;
        RECT  7.615 1.300 7.735 2.040 ;
        RECT  7.470 1.300 7.615 1.420 ;
        RECT  6.535 1.880 7.615 2.040 ;
        RECT  7.350 0.470 7.470 1.420 ;
        RECT  7.170 0.470 7.350 0.620 ;
        RECT  6.590 0.470 7.170 0.600 ;
        RECT  6.350 0.470 6.590 0.630 ;
        RECT  8.260 0.450 8.380 1.740 ;
        RECT  8.140 0.450 8.260 0.610 ;
        RECT  7.795 0.910 8.260 1.030 ;
        RECT  8.105 1.580 8.260 1.740 ;
        RECT  6.375 1.540 6.535 2.040 ;
        RECT  7.070 0.870 7.230 1.680 ;
        RECT  4.950 1.150 5.060 1.310 ;
        RECT  4.515 1.760 4.635 1.920 ;
        RECT  3.835 1.500 3.985 1.660 ;
        RECT  2.785 1.640 2.860 2.070 ;
        RECT  3.125 1.640 3.550 1.760 ;
        RECT  1.090 0.530 1.130 0.770 ;
        RECT  1.370 1.100 1.530 1.520 ;
        RECT  0.090 1.550 0.250 2.050 ;
        RECT  7.635 0.910 7.795 1.180 ;
        LAYER M1 ;
        RECT  8.810 0.490 9.015 0.870 ;
        RECT  8.790 1.650 9.015 2.030 ;
    END
END SDFKCNQD4

MACRO SDFKCSND1
    CLASS CORE ;
    FOREIGN SDFKCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.725 2.810 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.000 3.290 1.220 ;
        RECT  3.290 0.725 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.020 1.530 9.050 2.030 ;
        RECT  9.020 0.420 9.050 0.900 ;
        RECT  9.050 0.420 9.180 2.030 ;
        RECT  9.180 0.780 9.190 1.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.300 1.530 8.410 1.750 ;
        RECT  8.320 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.480 1.750 ;
        RECT  8.480 0.780 8.550 1.750 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.390 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.440 1.650 ;
        RECT  0.870 0.930 1.440 1.050 ;
        RECT  1.440 0.930 1.560 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.730 0.300 ;
        RECT  2.730 -0.300 2.950 0.490 ;
        RECT  2.950 -0.300 4.370 0.300 ;
        RECT  4.370 -0.300 4.590 0.350 ;
        RECT  4.590 -0.300 6.190 0.300 ;
        RECT  6.190 -0.300 6.410 0.760 ;
        RECT  6.410 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.740 2.820 ;
        RECT  2.740 2.030 2.960 2.820 ;
        RECT  2.960 2.220 3.345 2.820 ;
        RECT  3.345 2.160 3.565 2.820 ;
        RECT  3.565 2.220 4.415 2.820 ;
        RECT  4.415 2.160 4.635 2.820 ;
        RECT  4.635 2.220 6.125 2.820 ;
        RECT  6.125 1.760 6.345 2.820 ;
        RECT  6.345 2.220 7.555 2.820 ;
        RECT  7.555 2.160 7.775 2.820 ;
        RECT  7.775 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.885 1.580 8.040 1.740 ;
        RECT  7.575 0.910 8.040 1.030 ;
        RECT  7.920 0.450 8.040 0.610 ;
        RECT  8.040 0.450 8.160 2.050 ;
        RECT  8.160 1.930 8.715 2.050 ;
        RECT  8.715 1.050 8.835 2.050 ;
        RECT  8.835 1.050 8.930 1.270 ;
        RECT  7.120 0.460 7.240 1.420 ;
        RECT  6.865 1.880 7.395 2.040 ;
        RECT  7.240 1.300 7.395 1.420 ;
        RECT  7.395 1.300 7.515 2.040 ;
        RECT  7.515 1.300 7.735 1.420 ;
        RECT  7.735 1.160 7.895 1.420 ;
        RECT  7.000 1.540 7.100 1.680 ;
        RECT  7.100 1.540 7.255 1.760 ;
        RECT  6.020 1.150 6.150 1.580 ;
        RECT  6.150 1.460 6.535 1.580 ;
        RECT  6.535 1.460 6.590 1.980 ;
        RECT  6.590 0.540 6.710 1.980 ;
        RECT  6.710 0.540 6.760 0.780 ;
        RECT  5.580 0.590 5.595 0.830 ;
        RECT  5.595 0.590 5.715 1.920 ;
        RECT  5.715 0.590 5.740 1.020 ;
        RECT  5.740 0.900 6.300 1.020 ;
        RECT  6.300 0.900 6.460 1.300 ;
        RECT  4.750 0.740 4.945 0.900 ;
        RECT  4.945 0.740 5.065 1.660 ;
        RECT  5.065 1.130 5.465 1.290 ;
        RECT  3.690 0.430 3.820 0.850 ;
        RECT  3.820 0.430 3.910 2.070 ;
        RECT  3.910 0.470 3.945 2.070 ;
        RECT  3.945 1.640 3.965 2.070 ;
        RECT  3.965 1.890 5.095 2.010 ;
        RECT  3.945 0.470 5.170 0.590 ;
        RECT  5.095 1.890 5.335 2.050 ;
        RECT  5.170 0.450 5.410 0.620 ;
        RECT  4.080 0.720 4.510 0.880 ;
        RECT  4.510 0.720 4.630 1.760 ;
        RECT  4.630 1.050 4.795 1.270 ;
        RECT  2.210 0.600 2.330 0.760 ;
        RECT  2.210 1.730 3.415 1.890 ;
        RECT  3.415 1.370 3.535 1.890 ;
        RECT  3.535 1.370 3.550 1.490 ;
        RECT  3.550 0.970 3.690 1.490 ;
        RECT  2.490 1.365 2.930 1.520 ;
        RECT  2.930 0.660 3.050 1.520 ;
        RECT  3.050 0.660 3.170 0.880 ;
        RECT  3.050 1.360 3.280 1.520 ;
        RECT  1.240 1.930 1.740 2.050 ;
        RECT  1.040 0.620 1.740 0.780 ;
        RECT  1.740 0.420 1.900 2.050 ;
        RECT  0.060 0.590 0.350 0.750 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.320 1.310 ;
        RECT  6.930 0.460 7.120 0.620 ;
        RECT  6.840 0.870 7.000 1.680 ;
        RECT  5.910 1.150 6.020 1.310 ;
        RECT  5.475 1.760 5.595 1.920 ;
        RECT  4.795 1.500 4.945 1.660 ;
        RECT  3.745 1.640 3.820 2.070 ;
        RECT  4.085 1.640 4.510 1.760 ;
        RECT  2.090 0.600 2.210 1.890 ;
        RECT  2.330 1.100 2.490 1.520 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  0.070 1.850 0.350 2.010 ;
        RECT  7.415 0.910 7.575 1.180 ;
    END
END SDFKCSND1

MACRO SDFKCSND2
    CLASS CORE ;
    FOREIGN SDFKCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.725 2.810 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.000 3.290 1.220 ;
        RECT  3.290 0.725 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.280 1.950 9.310 2.090 ;
        RECT  9.310 1.380 9.370 2.090 ;
        RECT  9.310 0.420 9.370 0.900 ;
        RECT  9.370 0.420 9.470 2.090 ;
        RECT  9.470 1.950 9.500 2.090 ;
        RECT  9.470 0.780 9.510 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.410 8.730 1.570 ;
        RECT  8.610 0.420 8.730 0.900 ;
        RECT  8.730 0.420 8.770 1.570 ;
        RECT  8.770 0.780 8.870 1.570 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.390 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.500 1.650 ;
        RECT  0.870 0.930 1.500 1.050 ;
        RECT  1.500 0.930 1.620 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.730 0.300 ;
        RECT  2.730 -0.300 2.950 0.490 ;
        RECT  2.950 -0.300 4.370 0.300 ;
        RECT  4.370 -0.300 4.590 0.350 ;
        RECT  4.590 -0.300 6.190 0.300 ;
        RECT  6.190 -0.300 6.410 0.760 ;
        RECT  6.410 -0.300 9.920 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.740 2.820 ;
        RECT  2.740 2.030 2.960 2.820 ;
        RECT  2.960 2.220 3.345 2.820 ;
        RECT  3.345 2.160 3.565 2.820 ;
        RECT  3.565 2.220 4.415 2.820 ;
        RECT  4.415 2.160 4.635 2.820 ;
        RECT  4.635 2.220 6.125 2.820 ;
        RECT  6.125 1.760 6.345 2.820 ;
        RECT  6.345 2.220 7.555 2.820 ;
        RECT  7.555 2.160 7.775 2.820 ;
        RECT  7.775 2.220 8.160 2.820 ;
        RECT  8.160 2.160 8.380 2.820 ;
        RECT  8.380 2.220 9.920 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.590 0.540 6.710 1.980 ;
        RECT  6.710 0.540 6.760 0.780 ;
        RECT  5.580 0.590 5.595 0.830 ;
        RECT  5.595 0.590 5.715 1.920 ;
        RECT  5.715 0.590 5.740 1.020 ;
        RECT  5.740 0.900 6.300 1.020 ;
        RECT  6.300 0.900 6.460 1.300 ;
        RECT  4.750 0.740 4.945 0.900 ;
        RECT  4.945 0.740 5.065 1.660 ;
        RECT  5.065 1.130 5.465 1.290 ;
        RECT  3.690 0.430 3.820 0.850 ;
        RECT  3.820 0.430 3.910 2.070 ;
        RECT  3.910 0.470 3.945 2.070 ;
        RECT  3.945 1.640 3.965 2.070 ;
        RECT  3.965 1.890 5.095 2.010 ;
        RECT  3.945 0.470 5.170 0.590 ;
        RECT  5.095 1.890 5.335 2.050 ;
        RECT  5.170 0.450 5.410 0.620 ;
        RECT  4.080 0.720 4.510 0.880 ;
        RECT  4.510 0.720 4.630 1.760 ;
        RECT  4.630 1.050 4.795 1.270 ;
        RECT  2.210 0.600 2.330 0.760 ;
        RECT  2.210 1.730 3.415 1.890 ;
        RECT  3.415 1.370 3.535 1.890 ;
        RECT  3.535 1.370 3.550 1.490 ;
        RECT  3.550 0.970 3.690 1.490 ;
        RECT  2.490 1.365 2.930 1.520 ;
        RECT  2.930 0.660 3.050 1.520 ;
        RECT  3.050 0.660 3.170 0.880 ;
        RECT  3.050 1.360 3.280 1.520 ;
        RECT  1.240 1.930 1.740 2.050 ;
        RECT  1.040 0.620 1.740 0.780 ;
        RECT  1.740 0.420 1.900 2.050 ;
        RECT  0.060 0.590 0.350 0.750 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.380 1.310 ;
        RECT  6.535 1.460 6.590 1.980 ;
        RECT  6.150 1.460 6.535 1.580 ;
        RECT  6.020 1.150 6.150 1.580 ;
        RECT  7.100 1.540 7.255 1.760 ;
        RECT  7.000 1.540 7.100 1.680 ;
        RECT  7.735 1.160 7.895 1.420 ;
        RECT  7.515 1.300 7.735 1.420 ;
        RECT  7.395 1.300 7.515 2.040 ;
        RECT  7.240 1.300 7.395 1.420 ;
        RECT  6.865 1.880 7.395 2.040 ;
        RECT  7.120 0.460 7.240 1.420 ;
        RECT  9.125 1.050 9.220 1.270 ;
        RECT  9.005 1.050 9.125 1.810 ;
        RECT  8.160 1.690 9.005 1.810 ;
        RECT  8.040 0.450 8.160 1.810 ;
        RECT  7.890 0.450 8.040 0.610 ;
        RECT  7.575 0.910 8.040 1.030 ;
        RECT  7.885 1.580 8.040 1.740 ;
        RECT  6.930 0.460 7.120 0.620 ;
        RECT  6.840 0.870 7.000 1.680 ;
        RECT  5.910 1.150 6.020 1.310 ;
        RECT  5.475 1.760 5.595 1.920 ;
        RECT  4.795 1.500 4.945 1.660 ;
        RECT  3.745 1.640 3.820 2.070 ;
        RECT  4.085 1.640 4.510 1.760 ;
        RECT  2.090 0.600 2.210 1.890 ;
        RECT  2.330 1.100 2.490 1.520 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  0.070 1.850 0.350 2.010 ;
        RECT  7.415 0.910 7.575 1.180 ;
    END
END SDFKCSND2

MACRO SDFKCSND4
    CLASS CORE ;
    FOREIGN SDFKCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.230 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.650 0.725 2.810 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.000 3.290 1.220 ;
        RECT  3.290 0.725 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.130 1.650 11.470 2.030 ;
        RECT  11.150 0.490 11.470 0.870 ;
        RECT  11.470 0.490 11.890 2.030 ;
        RECT  11.890 1.650 12.060 2.030 ;
        RECT  11.890 0.490 12.060 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.730 1.560 9.870 1.720 ;
        RECT  9.770 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 1.720 ;
        RECT  10.290 1.560 10.680 1.720 ;
        RECT  10.290 0.490 10.680 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.565 0.890 1.795 ;
        RECT  0.890 1.490 1.110 1.795 ;
        RECT  1.110 1.565 1.190 1.795 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.250 1.005 4.390 1.515 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.590 0.890 0.730 1.130 ;
        RECT  0.730 0.445 0.870 1.050 ;
        RECT  1.320 1.490 1.500 1.650 ;
        RECT  0.870 0.930 1.500 1.050 ;
        RECT  1.500 0.930 1.620 1.650 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 2.730 0.300 ;
        RECT  2.730 -0.300 2.950 0.490 ;
        RECT  2.950 -0.300 6.190 0.300 ;
        RECT  6.190 -0.300 6.410 0.760 ;
        RECT  6.410 -0.300 6.970 0.300 ;
        RECT  6.970 -0.300 7.190 0.740 ;
        RECT  7.190 -0.300 12.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 2.790 2.820 ;
        RECT  2.790 2.030 3.010 2.820 ;
        RECT  3.010 2.220 3.345 2.820 ;
        RECT  3.345 2.160 3.565 2.820 ;
        RECT  3.565 2.220 6.125 2.820 ;
        RECT  6.125 1.760 6.345 2.820 ;
        RECT  6.345 2.220 6.885 2.820 ;
        RECT  6.885 1.760 7.105 2.820 ;
        RECT  7.105 2.220 8.735 2.820 ;
        RECT  8.735 2.160 8.955 2.820 ;
        RECT  8.955 2.220 9.350 2.820 ;
        RECT  9.350 2.160 9.570 2.820 ;
        RECT  9.570 2.220 12.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.910 0.470 3.945 2.070 ;
        RECT  3.945 1.640 3.965 2.070 ;
        RECT  3.965 1.890 5.095 2.010 ;
        RECT  3.945 0.470 5.170 0.590 ;
        RECT  5.095 1.890 5.335 2.050 ;
        RECT  5.170 0.470 5.410 0.630 ;
        RECT  4.080 0.720 4.510 0.880 ;
        RECT  4.510 0.720 4.630 1.760 ;
        RECT  4.630 1.050 4.795 1.270 ;
        RECT  2.210 0.600 2.330 0.760 ;
        RECT  2.210 1.730 3.415 1.890 ;
        RECT  3.415 1.370 3.535 1.890 ;
        RECT  3.535 1.370 3.550 1.490 ;
        RECT  3.550 0.970 3.690 1.490 ;
        RECT  2.490 1.365 2.930 1.520 ;
        RECT  2.930 0.660 3.050 1.520 ;
        RECT  3.050 0.660 3.170 0.880 ;
        RECT  3.050 1.360 3.280 1.520 ;
        RECT  1.240 1.930 1.740 2.050 ;
        RECT  1.040 0.620 1.740 0.780 ;
        RECT  1.740 0.420 1.900 2.050 ;
        RECT  0.060 0.590 0.350 0.750 ;
        RECT  0.350 0.590 0.470 2.010 ;
        RECT  0.470 1.280 0.640 1.440 ;
        RECT  0.640 1.250 0.760 1.440 ;
        RECT  0.760 1.250 0.950 1.370 ;
        RECT  0.950 1.170 1.070 1.370 ;
        RECT  1.070 1.170 1.380 1.310 ;
        RECT  3.820 0.430 3.910 2.070 ;
        RECT  3.690 0.430 3.820 0.850 ;
        RECT  5.065 1.130 5.465 1.290 ;
        RECT  4.945 0.740 5.065 1.660 ;
        RECT  4.750 0.740 4.945 0.900 ;
        RECT  6.300 0.900 6.460 1.300 ;
        RECT  5.740 0.900 6.300 1.020 ;
        RECT  5.715 0.590 5.740 1.020 ;
        RECT  5.595 0.590 5.715 1.920 ;
        RECT  5.580 0.590 5.595 0.830 ;
        RECT  7.875 0.720 7.900 0.940 ;
        RECT  7.760 0.720 7.875 1.760 ;
        RECT  7.715 0.860 7.760 1.760 ;
        RECT  6.760 0.860 7.715 0.980 ;
        RECT  6.710 0.540 6.760 0.980 ;
        RECT  6.590 0.540 6.710 1.980 ;
        RECT  6.535 1.460 6.590 1.980 ;
        RECT  6.150 1.460 6.535 1.580 ;
        RECT  6.020 1.150 6.150 1.580 ;
        RECT  8.280 1.540 8.435 1.760 ;
        RECT  8.190 1.540 8.280 1.680 ;
        RECT  8.915 1.160 9.075 1.420 ;
        RECT  8.695 1.300 8.915 1.420 ;
        RECT  8.575 1.300 8.695 2.040 ;
        RECT  8.430 1.300 8.575 1.420 ;
        RECT  7.495 1.880 8.575 2.040 ;
        RECT  8.310 0.470 8.430 1.420 ;
        RECT  8.130 0.470 8.310 0.620 ;
        RECT  7.550 0.470 8.130 0.600 ;
        RECT  7.310 0.470 7.550 0.630 ;
        RECT  11.005 1.050 11.190 1.270 ;
        RECT  10.885 1.050 11.005 2.040 ;
        RECT  9.340 1.920 10.885 2.040 ;
        RECT  9.220 0.450 9.340 2.040 ;
        RECT  9.100 0.450 9.220 0.610 ;
        RECT  8.755 0.910 9.220 1.030 ;
        RECT  9.065 1.580 9.220 1.740 ;
        RECT  7.335 1.540 7.495 2.040 ;
        RECT  8.030 0.870 8.190 1.680 ;
        RECT  5.910 1.150 6.020 1.310 ;
        RECT  5.475 1.760 5.595 1.920 ;
        RECT  4.795 1.500 4.945 1.660 ;
        RECT  3.745 1.640 3.820 2.070 ;
        RECT  4.085 1.640 4.510 1.760 ;
        RECT  2.090 0.600 2.210 1.890 ;
        RECT  8.595 0.910 8.755 1.180 ;
        RECT  2.330 1.110 2.490 1.520 ;
        RECT  1.000 1.930 1.240 2.090 ;
        RECT  0.070 1.850 0.350 2.010 ;
        LAYER M1 ;
        RECT  11.150 0.490 11.255 0.870 ;
        RECT  11.130 1.650 11.255 2.030 ;
        RECT  10.505 1.560 10.680 1.720 ;
        RECT  10.505 0.490 10.680 0.870 ;
    END
END SDFKCSND4

MACRO SDFKSND1
    CLASS CORE ;
    FOREIGN SDFKSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.285 0.550 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.725 2.490 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.020 2.970 1.180 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.670 1.940 8.700 2.100 ;
        RECT  8.700 1.390 8.730 2.100 ;
        RECT  8.700 0.440 8.730 0.940 ;
        RECT  8.730 0.440 8.860 2.100 ;
        RECT  8.860 0.820 8.870 1.515 ;
        RECT  8.860 1.940 8.890 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.960 1.550 8.090 1.770 ;
        RECT  7.980 0.420 8.090 0.920 ;
        RECT  8.090 0.420 8.140 1.770 ;
        RECT  8.140 0.800 8.230 1.770 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.345 ;
        RECT  0.570 -0.300 0.990 0.300 ;
        RECT  0.990 -0.300 1.210 0.345 ;
        RECT  1.210 -0.300 2.470 0.300 ;
        RECT  2.470 -0.300 2.690 0.490 ;
        RECT  2.690 -0.300 4.050 0.300 ;
        RECT  4.050 -0.300 4.270 0.340 ;
        RECT  4.270 -0.300 5.870 0.300 ;
        RECT  5.870 -0.300 6.090 0.760 ;
        RECT  6.090 -0.300 8.960 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.500 2.820 ;
        RECT  0.500 2.180 0.720 2.820 ;
        RECT  0.720 2.220 2.360 2.820 ;
        RECT  2.360 2.030 2.580 2.820 ;
        RECT  2.580 2.220 3.025 2.820 ;
        RECT  3.025 2.160 3.245 2.820 ;
        RECT  3.245 2.220 4.095 2.820 ;
        RECT  4.095 2.180 4.315 2.820 ;
        RECT  4.315 2.220 5.805 2.820 ;
        RECT  5.805 1.760 6.025 2.820 ;
        RECT  6.025 2.220 7.235 2.820 ;
        RECT  7.235 2.180 7.455 2.820 ;
        RECT  7.455 2.220 8.960 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.690 1.540 6.780 1.680 ;
        RECT  6.780 1.540 6.935 1.760 ;
        RECT  5.700 1.150 5.830 1.580 ;
        RECT  5.830 1.460 6.215 1.580 ;
        RECT  6.215 1.460 6.270 1.980 ;
        RECT  6.270 0.540 6.390 1.980 ;
        RECT  6.390 0.540 6.440 0.780 ;
        RECT  5.260 0.590 5.275 0.830 ;
        RECT  5.275 0.590 5.395 1.920 ;
        RECT  5.395 0.590 5.420 1.020 ;
        RECT  5.420 0.900 5.980 1.020 ;
        RECT  5.980 0.900 6.140 1.300 ;
        RECT  3.410 0.420 3.650 0.590 ;
        RECT  3.645 1.890 4.775 2.010 ;
        RECT  3.650 0.470 4.850 0.590 ;
        RECT  4.775 1.890 4.935 2.050 ;
        RECT  4.935 1.420 5.020 2.050 ;
        RECT  4.850 0.470 5.020 0.630 ;
        RECT  5.020 0.470 5.055 2.050 ;
        RECT  5.055 0.470 5.140 1.540 ;
        RECT  4.430 0.740 4.625 0.900 ;
        RECT  4.625 0.740 4.745 1.660 ;
        RECT  4.745 1.130 4.885 1.290 ;
        RECT  3.760 0.720 4.190 0.880 ;
        RECT  4.190 0.720 4.310 1.760 ;
        RECT  4.310 1.050 4.475 1.270 ;
        RECT  1.860 0.580 2.010 0.740 ;
        RECT  1.860 1.730 3.095 1.890 ;
        RECT  3.095 1.370 3.215 1.890 ;
        RECT  3.215 1.370 3.550 1.490 ;
        RECT  3.550 0.990 3.690 1.490 ;
        RECT  2.140 1.365 2.610 1.520 ;
        RECT  2.610 0.660 2.730 1.520 ;
        RECT  2.730 0.660 2.920 0.880 ;
        RECT  2.730 1.360 2.960 1.520 ;
        RECT  0.730 0.720 1.420 0.880 ;
        RECT  1.420 0.420 1.550 2.060 ;
        RECT  1.550 0.420 1.580 1.760 ;
        RECT  0.080 1.655 0.690 1.815 ;
        RECT  0.250 1.040 0.690 1.160 ;
        RECT  0.690 1.040 0.850 1.815 ;
        RECT  7.415 1.160 7.575 1.420 ;
        RECT  7.195 1.300 7.415 1.420 ;
        RECT  7.075 1.300 7.195 2.040 ;
        RECT  6.930 1.300 7.075 1.420 ;
        RECT  6.545 1.880 7.075 2.040 ;
        RECT  6.810 0.470 6.930 1.420 ;
        RECT  8.495 1.050 8.610 1.270 ;
        RECT  8.375 1.050 8.495 2.050 ;
        RECT  7.840 1.930 8.375 2.050 ;
        RECT  7.720 0.450 7.840 2.050 ;
        RECT  7.570 0.450 7.720 0.610 ;
        RECT  7.255 0.910 7.720 1.030 ;
        RECT  7.565 1.580 7.720 1.740 ;
        RECT  6.610 0.470 6.810 0.620 ;
        RECT  6.530 0.870 6.690 1.680 ;
        RECT  5.590 1.150 5.700 1.310 ;
        RECT  5.175 1.760 5.275 1.920 ;
        RECT  3.425 1.640 3.645 2.070 ;
        RECT  4.475 1.500 4.625 1.660 ;
        RECT  3.765 1.640 4.190 1.760 ;
        RECT  1.710 0.580 1.860 1.890 ;
        RECT  7.095 0.910 7.255 1.180 ;
        RECT  1.980 1.080 2.140 1.520 ;
        RECT  1.330 1.640 1.420 2.060 ;
        RECT  0.090 0.670 0.250 1.160 ;
    END
END SDFKSND1

MACRO SDFKSND2
    CLASS CORE ;
    FOREIGN SDFKSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.285 0.550 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.725 2.490 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.020 2.970 1.180 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.940 8.990 2.100 ;
        RECT  8.990 1.390 9.150 2.100 ;
        RECT  8.990 0.440 9.150 0.940 ;
        RECT  9.150 1.940 9.180 2.100 ;
        RECT  9.150 1.390 9.370 1.515 ;
        RECT  9.150 0.820 9.370 0.940 ;
        RECT  9.370 0.820 9.510 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.090 0.800 8.230 1.530 ;
        RECT  8.230 1.410 8.250 1.530 ;
        RECT  8.230 0.800 8.270 0.920 ;
        RECT  8.250 1.410 8.470 1.810 ;
        RECT  8.270 0.500 8.490 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.345 ;
        RECT  0.570 -0.300 0.990 0.300 ;
        RECT  0.990 -0.300 1.210 0.345 ;
        RECT  1.210 -0.300 2.470 0.300 ;
        RECT  2.470 -0.300 2.690 0.490 ;
        RECT  2.690 -0.300 4.050 0.300 ;
        RECT  4.050 -0.300 4.270 0.340 ;
        RECT  4.270 -0.300 5.870 0.300 ;
        RECT  5.870 -0.300 6.090 0.760 ;
        RECT  6.090 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.500 2.820 ;
        RECT  0.500 2.180 0.720 2.820 ;
        RECT  0.720 2.220 2.360 2.820 ;
        RECT  2.360 2.030 2.580 2.820 ;
        RECT  2.580 2.220 3.025 2.820 ;
        RECT  3.025 2.160 3.245 2.820 ;
        RECT  3.245 2.220 4.095 2.820 ;
        RECT  4.095 2.180 4.315 2.820 ;
        RECT  4.315 2.220 5.805 2.820 ;
        RECT  5.805 1.760 6.025 2.820 ;
        RECT  6.025 2.220 7.235 2.820 ;
        RECT  7.235 2.180 7.455 2.820 ;
        RECT  7.455 2.220 7.850 2.820 ;
        RECT  7.850 2.180 8.070 2.820 ;
        RECT  8.070 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.645 1.890 4.775 2.010 ;
        RECT  3.650 0.470 4.850 0.590 ;
        RECT  4.775 1.890 4.935 2.050 ;
        RECT  4.935 1.420 5.020 2.050 ;
        RECT  4.850 0.470 5.020 0.630 ;
        RECT  5.020 0.470 5.055 2.050 ;
        RECT  5.055 0.470 5.140 1.540 ;
        RECT  4.430 0.740 4.625 0.900 ;
        RECT  4.625 0.740 4.745 1.660 ;
        RECT  4.745 1.130 4.885 1.290 ;
        RECT  3.760 0.720 4.190 0.880 ;
        RECT  4.190 0.720 4.310 1.760 ;
        RECT  4.310 1.050 4.475 1.270 ;
        RECT  1.850 0.580 2.010 0.740 ;
        RECT  1.850 1.700 3.095 1.860 ;
        RECT  3.095 1.370 3.215 1.860 ;
        RECT  3.215 1.370 3.550 1.490 ;
        RECT  3.550 0.990 3.690 1.490 ;
        RECT  2.130 1.365 2.610 1.520 ;
        RECT  2.610 0.660 2.730 1.520 ;
        RECT  2.730 0.660 2.920 0.880 ;
        RECT  2.730 1.360 2.960 1.520 ;
        RECT  0.730 0.720 1.420 0.880 ;
        RECT  1.420 0.420 1.550 2.060 ;
        RECT  1.550 0.420 1.580 1.760 ;
        RECT  0.080 1.655 0.690 1.815 ;
        RECT  0.250 1.040 0.690 1.160 ;
        RECT  0.690 1.040 0.850 1.815 ;
        RECT  3.410 0.420 3.650 0.590 ;
        RECT  5.980 0.900 6.140 1.300 ;
        RECT  5.420 0.900 5.980 1.020 ;
        RECT  5.395 0.590 5.420 1.020 ;
        RECT  5.275 0.590 5.395 1.920 ;
        RECT  5.260 0.590 5.275 0.830 ;
        RECT  6.390 0.540 6.440 0.780 ;
        RECT  6.270 0.540 6.390 1.980 ;
        RECT  6.215 1.460 6.270 1.980 ;
        RECT  5.830 1.460 6.215 1.580 ;
        RECT  5.700 1.150 5.830 1.580 ;
        RECT  6.780 1.540 6.935 1.760 ;
        RECT  6.690 1.540 6.780 1.680 ;
        RECT  7.415 1.160 7.575 1.420 ;
        RECT  7.195 1.300 7.415 1.420 ;
        RECT  7.075 1.300 7.195 2.040 ;
        RECT  6.930 1.300 7.075 1.420 ;
        RECT  6.545 1.880 7.075 2.040 ;
        RECT  6.810 0.470 6.930 1.420 ;
        RECT  8.815 1.080 9.050 1.240 ;
        RECT  8.695 1.080 8.815 2.050 ;
        RECT  7.840 1.930 8.695 2.050 ;
        RECT  7.720 0.450 7.840 2.050 ;
        RECT  7.600 0.450 7.720 0.610 ;
        RECT  7.255 0.910 7.720 1.030 ;
        RECT  7.565 1.580 7.720 1.740 ;
        RECT  6.610 0.470 6.810 0.620 ;
        RECT  6.530 0.870 6.690 1.680 ;
        RECT  5.590 1.150 5.700 1.310 ;
        RECT  5.175 1.760 5.275 1.920 ;
        RECT  3.425 1.640 3.645 2.070 ;
        RECT  4.475 1.500 4.625 1.660 ;
        RECT  3.765 1.640 4.190 1.760 ;
        RECT  1.710 0.580 1.850 1.860 ;
        RECT  1.970 1.080 2.130 1.520 ;
        RECT  1.330 1.640 1.420 2.060 ;
        RECT  0.090 0.670 0.250 1.160 ;
        RECT  7.095 0.910 7.255 1.180 ;
    END
END SDFKSND2

MACRO SDFKSND4
    CLASS CORE ;
    FOREIGN SDFKSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.285 0.550 1.515 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 0.725 2.490 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.850 1.020 2.970 1.180 ;
        RECT  2.970 1.005 3.430 1.235 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.810 1.650 11.150 2.030 ;
        RECT  10.830 0.490 11.150 0.870 ;
        RECT  11.150 0.490 11.570 2.030 ;
        RECT  11.570 1.650 11.740 2.030 ;
        RECT  11.570 0.490 11.740 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.410 1.560 9.550 1.720 ;
        RECT  9.450 0.490 9.550 0.870 ;
        RECT  9.550 0.490 9.970 1.720 ;
        RECT  9.970 1.560 10.360 1.720 ;
        RECT  9.970 0.490 10.360 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.210 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.350 0.300 ;
        RECT  0.350 -0.300 0.570 0.345 ;
        RECT  0.570 -0.300 0.990 0.300 ;
        RECT  0.990 -0.300 1.210 0.345 ;
        RECT  1.210 -0.300 2.470 0.300 ;
        RECT  2.470 -0.300 2.690 0.490 ;
        RECT  2.690 -0.300 5.870 0.300 ;
        RECT  5.870 -0.300 6.090 0.760 ;
        RECT  6.090 -0.300 6.650 0.300 ;
        RECT  6.650 -0.300 6.870 0.740 ;
        RECT  6.870 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.500 2.820 ;
        RECT  0.500 2.180 0.720 2.820 ;
        RECT  0.720 2.220 2.360 2.820 ;
        RECT  2.360 2.030 2.580 2.820 ;
        RECT  2.580 2.220 3.025 2.820 ;
        RECT  3.025 2.160 3.245 2.820 ;
        RECT  3.245 2.220 5.805 2.820 ;
        RECT  5.805 1.760 6.025 2.820 ;
        RECT  6.025 2.220 6.565 2.820 ;
        RECT  6.565 1.760 6.785 2.820 ;
        RECT  6.785 2.220 8.415 2.820 ;
        RECT  8.415 2.160 8.635 2.820 ;
        RECT  8.635 2.220 9.030 2.820 ;
        RECT  9.030 2.160 9.250 2.820 ;
        RECT  9.250 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.690 1.040 0.850 1.815 ;
        RECT  0.250 1.040 0.690 1.160 ;
        RECT  0.080 1.655 0.690 1.815 ;
        RECT  1.550 0.420 1.580 1.760 ;
        RECT  1.420 0.420 1.550 2.060 ;
        RECT  0.730 0.720 1.420 0.880 ;
        RECT  2.730 1.360 2.960 1.520 ;
        RECT  2.730 0.660 2.920 0.880 ;
        RECT  2.610 0.660 2.730 1.520 ;
        RECT  2.130 1.365 2.610 1.520 ;
        RECT  3.550 0.990 3.690 1.490 ;
        RECT  3.215 1.370 3.550 1.490 ;
        RECT  3.095 1.370 3.215 1.860 ;
        RECT  1.850 1.700 3.095 1.860 ;
        RECT  1.850 0.580 2.010 0.740 ;
        RECT  4.310 1.050 4.475 1.270 ;
        RECT  4.190 0.720 4.310 1.760 ;
        RECT  3.760 0.720 4.190 0.880 ;
        RECT  4.745 1.130 4.885 1.290 ;
        RECT  4.625 0.740 4.745 1.660 ;
        RECT  4.430 0.740 4.625 0.900 ;
        RECT  5.055 0.470 5.140 1.540 ;
        RECT  5.020 0.470 5.055 2.050 ;
        RECT  4.850 0.470 5.020 0.630 ;
        RECT  4.935 1.420 5.020 2.050 ;
        RECT  4.775 1.890 4.935 2.050 ;
        RECT  3.650 0.470 4.850 0.590 ;
        RECT  3.645 1.890 4.775 2.010 ;
        RECT  3.410 0.420 3.650 0.590 ;
        RECT  5.980 0.900 6.140 1.300 ;
        RECT  5.420 0.900 5.980 1.020 ;
        RECT  5.395 0.590 5.420 1.020 ;
        RECT  5.275 0.590 5.395 1.920 ;
        RECT  5.260 0.590 5.275 0.830 ;
        RECT  7.555 0.720 7.580 0.940 ;
        RECT  7.440 0.720 7.555 1.760 ;
        RECT  7.395 0.860 7.440 1.760 ;
        RECT  6.440 0.860 7.395 0.980 ;
        RECT  6.390 0.540 6.440 0.980 ;
        RECT  6.270 0.540 6.390 1.980 ;
        RECT  6.215 1.460 6.270 1.980 ;
        RECT  5.830 1.460 6.215 1.580 ;
        RECT  5.700 1.150 5.830 1.580 ;
        RECT  7.960 1.540 8.115 1.760 ;
        RECT  7.870 1.540 7.960 1.680 ;
        RECT  8.595 1.160 8.755 1.420 ;
        RECT  8.375 1.300 8.595 1.420 ;
        RECT  8.255 1.300 8.375 2.040 ;
        RECT  8.110 1.300 8.255 1.420 ;
        RECT  7.175 1.880 8.255 2.040 ;
        RECT  7.990 0.470 8.110 1.420 ;
        RECT  7.810 0.470 7.990 0.620 ;
        RECT  7.230 0.470 7.810 0.600 ;
        RECT  6.990 0.470 7.230 0.630 ;
        RECT  10.685 1.050 10.870 1.270 ;
        RECT  10.565 1.050 10.685 2.040 ;
        RECT  9.020 1.920 10.565 2.040 ;
        RECT  8.900 0.450 9.020 2.040 ;
        RECT  8.780 0.450 8.900 0.610 ;
        RECT  8.435 0.910 8.900 1.030 ;
        RECT  8.745 1.580 8.900 1.740 ;
        RECT  7.015 1.540 7.175 2.040 ;
        RECT  7.710 0.870 7.870 1.680 ;
        RECT  5.590 1.150 5.700 1.310 ;
        RECT  5.175 1.760 5.275 1.920 ;
        RECT  3.425 1.640 3.645 2.070 ;
        RECT  4.475 1.500 4.625 1.660 ;
        RECT  3.765 1.640 4.190 1.760 ;
        RECT  1.710 0.580 1.850 1.860 ;
        RECT  1.970 1.080 2.130 1.520 ;
        RECT  1.330 1.640 1.420 2.060 ;
        RECT  0.090 0.670 0.250 1.160 ;
        RECT  8.275 0.910 8.435 1.180 ;
        LAYER M1 ;
        RECT  10.810 1.650 10.935 2.030 ;
        RECT  10.185 1.560 10.360 1.720 ;
        RECT  10.185 0.490 10.360 0.870 ;
        RECT  10.830 0.490 10.935 0.870 ;
    END
END SDFKSND4

MACRO SDFNCND1
    CLASS CORE ;
    FOREIGN SDFNCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.940 1.940 8.970 2.100 ;
        RECT  8.970 1.390 9.050 2.100 ;
        RECT  8.970 0.420 9.050 0.900 ;
        RECT  9.050 0.420 9.130 2.100 ;
        RECT  9.130 1.940 9.160 2.100 ;
        RECT  9.130 0.760 9.190 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.220 1.960 8.250 2.100 ;
        RECT  8.250 1.390 8.410 2.100 ;
        RECT  8.200 0.710 8.410 0.870 ;
        RECT  8.410 1.960 8.440 2.100 ;
        RECT  8.410 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.760 1.285 7.920 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.460 0.300 ;
        RECT  4.460 -0.300 4.610 0.720 ;
        RECT  4.610 -0.300 6.500 0.300 ;
        RECT  6.500 -0.300 6.720 0.590 ;
        RECT  6.720 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.940 2.820 ;
        RECT  4.940 2.040 5.160 2.820 ;
        RECT  5.160 2.220 6.500 2.820 ;
        RECT  6.500 2.180 6.720 2.820 ;
        RECT  6.720 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.810 1.650 7.110 1.810 ;
        RECT  6.810 0.950 7.140 1.070 ;
        RECT  7.140 0.710 7.360 1.070 ;
        RECT  7.360 0.950 7.480 1.070 ;
        RECT  7.480 0.950 7.600 2.050 ;
        RECT  7.600 1.930 7.820 2.050 ;
        RECT  7.600 1.020 8.070 1.160 ;
        RECT  8.070 1.020 8.290 1.180 ;
        RECT  5.510 1.190 5.750 1.310 ;
        RECT  5.750 1.190 5.910 2.050 ;
        RECT  5.910 1.930 7.230 2.050 ;
        RECT  7.190 1.290 7.230 1.530 ;
        RECT  7.230 1.290 7.350 2.050 ;
        RECT  3.850 0.430 3.970 0.960 ;
        RECT  3.970 0.840 4.730 0.960 ;
        RECT  4.730 0.470 4.850 0.960 ;
        RECT  4.850 0.470 5.810 0.610 ;
        RECT  5.810 0.450 6.030 0.610 ;
        RECT  4.310 1.420 5.090 1.580 ;
        RECT  4.970 0.730 5.090 0.950 ;
        RECT  5.090 0.730 5.230 1.580 ;
        RECT  5.230 1.440 5.370 1.580 ;
        RECT  5.370 1.440 5.530 1.960 ;
        RECT  3.610 0.710 3.720 1.910 ;
        RECT  3.720 1.080 3.770 1.910 ;
        RECT  3.770 1.080 4.830 1.200 ;
        RECT  4.830 1.080 4.970 1.300 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.100 3.430 1.260 ;
        RECT  1.410 1.930 3.190 2.050 ;
        RECT  3.190 1.930 3.430 2.090 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.510 0.710 1.630 0.870 ;
        RECT  1.630 0.710 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  6.670 0.950 6.810 1.810 ;
        RECT  8.850 1.050 8.890 1.290 ;
        RECT  8.710 0.470 8.850 1.290 ;
        RECT  7.000 0.470 8.710 0.590 ;
        RECT  6.880 0.470 7.000 0.830 ;
        RECT  6.330 0.710 6.880 0.830 ;
        RECT  6.170 0.650 6.330 0.975 ;
        RECT  6.170 1.510 6.270 1.730 ;
        RECT  6.160 0.650 6.170 1.730 ;
        RECT  6.030 0.820 6.160 1.730 ;
        RECT  5.680 0.820 6.030 0.980 ;
        RECT  6.310 1.125 6.670 1.345 ;
        RECT  5.350 0.770 5.510 1.310 ;
        RECT  3.700 0.430 3.850 0.590 ;
        RECT  4.090 1.410 4.310 1.580 ;
        RECT  3.560 0.710 3.610 1.195 ;
        RECT  3.940 1.700 4.910 1.860 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
    END
END SDFNCND1

MACRO SDFNCND2
    CLASS CORE ;
    FOREIGN SDFNCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.950 8.990 2.090 ;
        RECT  8.990 1.380 9.150 2.090 ;
        RECT  9.150 1.950 9.180 2.090 ;
        RECT  8.960 0.490 9.180 0.910 ;
        RECT  9.150 1.380 9.370 1.515 ;
        RECT  9.180 0.790 9.370 0.910 ;
        RECT  9.370 0.790 9.510 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.270 1.950 8.300 2.090 ;
        RECT  8.300 1.380 8.410 2.090 ;
        RECT  8.240 0.710 8.410 0.870 ;
        RECT  8.410 0.710 8.460 2.090 ;
        RECT  8.460 1.950 8.490 2.090 ;
        RECT  8.460 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.285 7.910 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.460 0.300 ;
        RECT  2.460 -0.300 2.680 0.340 ;
        RECT  2.680 -0.300 4.460 0.300 ;
        RECT  4.460 -0.300 4.610 0.720 ;
        RECT  4.610 -0.300 6.500 0.300 ;
        RECT  6.500 -0.300 6.720 0.590 ;
        RECT  6.720 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 2.000 2.820 ;
        RECT  2.000 2.180 2.220 2.820 ;
        RECT  2.220 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.940 2.820 ;
        RECT  4.940 2.040 5.160 2.820 ;
        RECT  5.160 2.220 6.500 2.820 ;
        RECT  6.500 2.180 6.720 2.820 ;
        RECT  6.720 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.120 1.020 8.290 1.180 ;
        RECT  5.510 1.190 5.750 1.310 ;
        RECT  5.750 1.190 5.910 2.050 ;
        RECT  5.910 1.930 7.230 2.050 ;
        RECT  7.190 1.290 7.230 1.530 ;
        RECT  7.230 1.290 7.350 2.050 ;
        RECT  3.850 0.430 3.970 0.960 ;
        RECT  3.970 0.840 4.730 0.960 ;
        RECT  4.730 0.470 4.850 0.960 ;
        RECT  4.850 0.470 5.810 0.610 ;
        RECT  5.810 0.450 6.030 0.610 ;
        RECT  4.310 1.420 5.090 1.580 ;
        RECT  4.970 0.730 5.090 0.950 ;
        RECT  5.090 0.730 5.230 1.580 ;
        RECT  5.230 1.440 5.370 1.580 ;
        RECT  5.370 1.440 5.530 1.960 ;
        RECT  3.610 0.710 3.720 1.910 ;
        RECT  3.720 1.080 3.770 1.910 ;
        RECT  3.770 1.080 4.830 1.200 ;
        RECT  4.830 1.080 4.970 1.300 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.100 3.430 1.260 ;
        RECT  1.410 1.930 3.190 2.050 ;
        RECT  3.190 1.930 3.430 2.090 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.710 1.630 0.870 ;
        RECT  1.630 0.710 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  8.000 0.710 8.120 1.180 ;
        RECT  7.600 0.710 8.000 0.830 ;
        RECT  7.600 1.930 7.820 2.050 ;
        RECT  7.480 0.710 7.600 2.050 ;
        RECT  7.170 0.710 7.480 1.070 ;
        RECT  6.810 0.950 7.170 1.070 ;
        RECT  6.810 1.650 7.110 1.810 ;
        RECT  6.670 0.950 6.810 1.810 ;
        RECT  8.840 1.080 9.080 1.240 ;
        RECT  8.720 0.470 8.840 1.240 ;
        RECT  7.000 0.470 8.720 0.590 ;
        RECT  6.880 0.470 7.000 0.830 ;
        RECT  6.330 0.710 6.880 0.830 ;
        RECT  6.170 0.650 6.330 0.975 ;
        RECT  6.170 1.510 6.270 1.730 ;
        RECT  6.160 0.650 6.170 1.730 ;
        RECT  6.030 0.820 6.160 1.730 ;
        RECT  6.310 1.125 6.670 1.345 ;
        RECT  5.350 0.770 5.510 1.310 ;
        RECT  5.680 0.820 6.030 0.980 ;
        RECT  3.690 0.430 3.850 0.590 ;
        RECT  4.090 1.410 4.310 1.580 ;
        RECT  3.560 0.710 3.610 1.195 ;
        RECT  3.940 1.700 4.910 1.860 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
    END
END SDFNCND2

MACRO SDFNCND4
    CLASS CORE ;
    FOREIGN SDFNCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.200 0.870 1.795 ;
        RECT  0.870 1.200 0.930 1.420 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 1.650 10.830 2.030 ;
        RECT  10.430 0.490 10.830 0.870 ;
        RECT  10.830 0.490 11.250 2.030 ;
        RECT  11.250 1.650 11.360 2.030 ;
        RECT  11.250 0.490 11.360 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.990 1.610 9.230 1.770 ;
        RECT  8.960 0.760 9.230 0.920 ;
        RECT  9.230 0.760 9.650 1.770 ;
        RECT  9.650 1.610 9.960 1.770 ;
        RECT  9.650 0.760 9.960 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.870 1.200 2.010 1.420 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.170 2.490 1.390 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.770 1.190 7.950 1.515 ;
        RECT  7.950 1.285 8.230 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.490 ;
        RECT  0.680 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.620 0.720 ;
        RECT  4.620 -0.300 6.510 0.300 ;
        RECT  6.510 -0.300 6.730 0.590 ;
        RECT  6.730 -0.300 7.790 0.300 ;
        RECT  7.790 -0.300 8.010 0.340 ;
        RECT  8.010 -0.300 8.590 0.300 ;
        RECT  8.590 -0.300 8.810 0.340 ;
        RECT  8.810 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 4.950 2.820 ;
        RECT  4.950 2.040 5.170 2.820 ;
        RECT  5.170 2.220 6.510 2.820 ;
        RECT  6.510 2.180 6.730 2.820 ;
        RECT  6.730 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.070 0.830 3.190 1.720 ;
        RECT  3.190 1.100 3.440 1.260 ;
        RECT  1.410 1.930 3.200 2.050 ;
        RECT  3.200 1.930 3.440 2.090 ;
        RECT  1.340 0.470 3.130 0.590 ;
        RECT  3.130 0.470 3.370 0.630 ;
        RECT  2.150 0.710 2.630 0.870 ;
        RECT  2.630 0.710 2.750 1.810 ;
        RECT  2.750 1.170 2.950 1.330 ;
        RECT  1.480 0.710 1.630 0.870 ;
        RECT  1.630 0.710 1.750 1.780 ;
        RECT  1.750 1.620 1.840 1.780 ;
        RECT  0.060 1.690 0.370 1.850 ;
        RECT  0.250 0.765 0.370 0.885 ;
        RECT  0.370 0.765 0.490 1.850 ;
        RECT  0.490 0.765 1.100 0.885 ;
        RECT  1.100 0.765 1.260 1.440 ;
        RECT  2.870 0.830 3.070 0.990 ;
        RECT  4.830 1.080 4.970 1.300 ;
        RECT  3.780 1.080 4.830 1.200 ;
        RECT  3.720 1.080 3.780 1.910 ;
        RECT  3.620 0.710 3.720 1.910 ;
        RECT  5.380 1.440 5.540 1.960 ;
        RECT  5.240 1.440 5.380 1.580 ;
        RECT  5.120 0.730 5.240 1.580 ;
        RECT  4.980 0.730 5.120 0.950 ;
        RECT  4.320 1.420 5.120 1.580 ;
        RECT  5.820 0.450 6.040 0.610 ;
        RECT  4.860 0.470 5.820 0.610 ;
        RECT  4.740 0.470 4.860 0.960 ;
        RECT  3.980 0.840 4.740 0.960 ;
        RECT  3.860 0.430 3.980 0.960 ;
        RECT  7.250 1.190 7.370 2.050 ;
        RECT  7.210 1.190 7.250 1.410 ;
        RECT  5.920 1.930 7.250 2.050 ;
        RECT  5.760 1.190 5.920 2.050 ;
        RECT  5.520 1.190 5.760 1.310 ;
        RECT  8.560 1.080 8.740 1.240 ;
        RECT  8.440 0.950 8.560 1.240 ;
        RECT  7.610 0.950 8.440 1.070 ;
        RECT  7.610 1.890 7.840 2.050 ;
        RECT  7.490 0.950 7.610 2.050 ;
        RECT  7.340 0.950 7.490 1.070 ;
        RECT  7.180 0.710 7.340 1.070 ;
        RECT  6.820 0.950 7.180 1.070 ;
        RECT  6.820 1.650 7.130 1.810 ;
        RECT  6.680 0.950 6.820 1.810 ;
        RECT  10.260 1.080 10.540 1.240 ;
        RECT  10.140 0.470 10.260 2.050 ;
        RECT  7.010 0.470 10.140 0.590 ;
        RECT  8.220 1.890 10.140 2.050 ;
        RECT  6.890 0.470 7.010 0.830 ;
        RECT  6.340 0.710 6.890 0.830 ;
        RECT  6.180 0.650 6.340 0.975 ;
        RECT  6.180 1.495 6.280 1.715 ;
        RECT  6.170 0.650 6.180 1.715 ;
        RECT  6.040 0.820 6.170 1.715 ;
        RECT  6.320 1.125 6.680 1.345 ;
        RECT  5.690 0.820 6.040 0.980 ;
        RECT  5.360 0.770 5.520 1.310 ;
        RECT  3.710 0.430 3.860 0.590 ;
        RECT  4.100 1.410 4.320 1.580 ;
        RECT  3.560 0.710 3.620 1.195 ;
        RECT  3.950 1.700 4.920 1.860 ;
        RECT  2.910 1.560 3.070 1.720 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.100 0.430 1.340 0.590 ;
        RECT  2.220 1.650 2.630 1.810 ;
        RECT  1.600 1.620 1.630 1.780 ;
        RECT  0.090 0.570 0.250 0.885 ;
        LAYER M1 ;
        RECT  10.430 1.650 10.615 2.030 ;
        RECT  10.430 0.490 10.615 0.870 ;
        RECT  9.865 1.610 9.960 1.770 ;
        RECT  9.865 0.760 9.960 0.920 ;
        RECT  8.990 1.610 9.015 1.770 ;
        RECT  8.960 0.760 9.015 0.920 ;
    END
END SDFNCND4

MACRO SDFNCSND1
    CLASS CORE ;
    FOREIGN SDFNCSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.080 0.725 8.240 1.290 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.600 1.490 8.730 1.650 ;
        RECT  8.630 0.420 8.730 0.910 ;
        RECT  8.730 0.420 8.790 1.650 ;
        RECT  8.790 0.790 8.870 1.650 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.320 1.960 9.350 2.100 ;
        RECT  9.350 1.390 9.370 2.100 ;
        RECT  9.350 0.420 9.370 0.900 ;
        RECT  9.370 0.420 9.510 2.100 ;
        RECT  9.510 1.960 9.540 2.100 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 7.270 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 7.480 0.300 ;
        RECT  7.480 -0.300 7.700 0.340 ;
        RECT  7.700 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.470 2.820 ;
        RECT  2.470 2.180 2.690 2.820 ;
        RECT  2.690 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.760 2.820 ;
        RECT  6.760 1.970 6.980 2.820 ;
        RECT  6.980 2.220 7.560 2.820 ;
        RECT  7.560 2.010 7.780 2.820 ;
        RECT  7.780 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.580 1.450 6.750 1.610 ;
        RECT  6.580 0.470 8.250 0.590 ;
        RECT  7.940 1.490 8.360 1.650 ;
        RECT  8.250 0.430 8.360 0.590 ;
        RECT  8.360 0.430 8.480 1.650 ;
        RECT  8.480 1.050 8.610 1.270 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  6.220 1.160 6.340 2.040 ;
        RECT  6.340 1.730 6.440 2.040 ;
        RECT  6.440 1.730 6.870 1.850 ;
        RECT  6.870 1.490 6.990 1.850 ;
        RECT  6.990 1.490 7.390 1.610 ;
        RECT  7.390 1.030 7.550 1.610 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.940 1.780 6.100 2.090 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.050 3.240 1.270 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  6.460 0.470 6.580 1.610 ;
        RECT  9.220 1.030 9.250 1.270 ;
        RECT  9.100 1.030 9.220 1.890 ;
        RECT  7.790 1.770 9.100 1.890 ;
        RECT  7.790 1.080 7.960 1.240 ;
        RECT  7.670 0.710 7.790 1.890 ;
        RECT  6.790 0.710 7.670 0.870 ;
        RECT  7.140 1.730 7.670 1.890 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  3.690 1.930 3.930 2.090 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFNCSND1

MACRO SDFNCSND2
    CLASS CORE ;
    FOREIGN SDFNCSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.730 1.005 9.190 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.550 1.410 9.690 1.810 ;
        RECT  9.580 0.420 9.690 0.900 ;
        RECT  9.690 0.420 9.740 1.810 ;
        RECT  9.740 0.780 9.770 1.810 ;
        RECT  9.770 0.780 9.830 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.240 1.940 10.270 2.100 ;
        RECT  10.270 1.390 10.330 2.100 ;
        RECT  10.270 0.420 10.330 0.900 ;
        RECT  10.330 0.420 10.430 2.100 ;
        RECT  10.430 1.940 10.460 2.100 ;
        RECT  10.430 0.780 10.470 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.005 7.910 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.530 0.300 ;
        RECT  2.530 -0.300 2.750 0.340 ;
        RECT  2.750 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 6.970 0.300 ;
        RECT  6.970 -0.300 7.190 0.490 ;
        RECT  7.190 -0.300 8.260 0.300 ;
        RECT  8.260 -0.300 8.480 0.340 ;
        RECT  8.480 -0.300 9.150 0.300 ;
        RECT  9.150 -0.300 9.370 0.340 ;
        RECT  9.370 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.470 2.820 ;
        RECT  2.470 2.180 2.690 2.820 ;
        RECT  2.690 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.850 2.820 ;
        RECT  6.850 2.030 7.070 2.820 ;
        RECT  7.070 2.220 8.330 2.820 ;
        RECT  8.330 2.010 8.550 2.820 ;
        RECT  8.550 2.220 9.140 2.820 ;
        RECT  9.140 2.180 9.360 2.820 ;
        RECT  9.360 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.050 3.250 1.270 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  5.940 1.780 6.100 2.100 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  8.120 1.030 8.280 1.500 ;
        RECT  7.310 1.380 8.120 1.500 ;
        RECT  7.150 1.030 7.310 1.500 ;
        RECT  7.070 1.380 7.150 1.500 ;
        RECT  6.950 1.380 7.070 1.850 ;
        RECT  6.440 1.730 6.950 1.850 ;
        RECT  6.340 1.730 6.440 2.040 ;
        RECT  6.220 1.160 6.340 2.040 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  9.430 1.080 9.570 1.240 ;
        RECT  9.310 0.720 9.430 1.650 ;
        RECT  9.090 0.720 9.310 0.840 ;
        RECT  8.700 1.490 9.310 1.650 ;
        RECT  8.930 0.470 9.090 0.840 ;
        RECT  7.500 0.470 8.930 0.590 ;
        RECT  7.380 0.470 7.500 0.830 ;
        RECT  6.580 0.710 7.380 0.830 ;
        RECT  6.580 1.450 6.750 1.610 ;
        RECT  6.460 0.710 6.580 1.610 ;
        RECT  10.120 1.050 10.210 1.270 ;
        RECT  10.000 1.050 10.120 2.050 ;
        RECT  9.220 1.930 10.000 2.050 ;
        RECT  9.100 1.770 9.220 2.050 ;
        RECT  8.580 1.770 9.100 1.890 ;
        RECT  8.580 1.050 8.610 1.270 ;
        RECT  8.460 0.710 8.580 1.890 ;
        RECT  7.620 0.710 8.460 0.850 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  3.690 1.930 3.930 2.090 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  7.230 1.620 8.460 1.780 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFNCSND2

MACRO SDFNCSND4
    CLASS CORE ;
    FOREIGN SDFNCSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.730 0.725 8.870 1.235 ;
        RECT  8.870 1.075 9.005 1.235 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.430 1.600 9.870 1.760 ;
        RECT  9.450 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 1.760 ;
        RECT  10.290 0.490 10.360 0.870 ;
        RECT  10.290 1.600 10.380 1.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.830 1.650 11.150 2.030 ;
        RECT  10.830 0.490 11.150 0.870 ;
        RECT  11.150 0.490 11.570 2.030 ;
        RECT  11.570 1.650 11.740 2.030 ;
        RECT  11.570 0.490 11.740 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.450 1.005 7.910 1.235 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 4.760 0.300 ;
        RECT  4.760 -0.300 4.980 0.490 ;
        RECT  4.980 -0.300 6.880 0.300 ;
        RECT  6.880 -0.300 7.100 0.490 ;
        RECT  7.100 -0.300 8.170 0.300 ;
        RECT  8.170 -0.300 8.390 0.340 ;
        RECT  8.390 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 4.780 2.820 ;
        RECT  4.780 2.180 5.000 2.820 ;
        RECT  5.000 2.220 5.580 2.820 ;
        RECT  5.580 2.020 5.800 2.820 ;
        RECT  5.800 2.220 6.760 2.820 ;
        RECT  6.760 2.030 6.980 2.820 ;
        RECT  6.980 2.220 8.240 2.820 ;
        RECT  8.240 2.010 8.460 2.820 ;
        RECT  8.460 2.220 9.040 2.820 ;
        RECT  9.040 2.180 9.260 2.820 ;
        RECT  9.260 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.680 1.500 6.060 1.660 ;
        RECT  4.030 0.430 4.150 0.730 ;
        RECT  4.150 0.610 5.100 0.730 ;
        RECT  5.100 0.470 5.220 0.730 ;
        RECT  5.220 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  3.630 1.040 3.720 1.810 ;
        RECT  3.720 0.720 3.750 1.810 ;
        RECT  3.750 0.720 3.880 1.180 ;
        RECT  3.880 1.040 5.230 1.180 ;
        RECT  4.420 1.540 4.540 1.810 ;
        RECT  4.540 1.540 4.710 1.700 ;
        RECT  1.380 0.470 3.330 0.590 ;
        RECT  3.330 0.470 3.490 0.840 ;
        RECT  1.280 1.920 3.130 2.040 ;
        RECT  3.130 1.920 3.370 2.080 ;
        RECT  2.920 0.710 3.050 0.870 ;
        RECT  3.050 0.710 3.170 1.660 ;
        RECT  3.170 1.030 3.270 1.250 ;
        RECT  2.230 0.710 2.610 0.870 ;
        RECT  2.610 0.710 2.730 1.800 ;
        RECT  2.730 1.050 2.920 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  5.520 0.710 5.680 1.660 ;
        RECT  4.980 1.500 5.520 1.660 ;
        RECT  4.860 1.300 4.980 1.660 ;
        RECT  4.330 1.300 4.860 1.420 ;
        RECT  5.940 1.780 6.100 2.100 ;
        RECT  5.320 1.780 5.940 1.900 ;
        RECT  5.200 1.780 5.320 2.050 ;
        RECT  3.930 1.930 5.200 2.050 ;
        RECT  8.030 1.030 8.190 1.500 ;
        RECT  7.220 1.380 8.030 1.500 ;
        RECT  7.060 1.030 7.220 1.500 ;
        RECT  6.980 1.380 7.060 1.500 ;
        RECT  6.860 1.380 6.980 1.850 ;
        RECT  6.440 1.730 6.860 1.850 ;
        RECT  6.340 1.730 6.440 2.040 ;
        RECT  6.220 1.160 6.340 2.040 ;
        RECT  6.060 1.160 6.220 1.280 ;
        RECT  9.245 1.080 9.570 1.240 ;
        RECT  9.125 0.430 9.245 1.650 ;
        RECT  8.810 0.430 9.125 0.590 ;
        RECT  8.610 1.490 9.125 1.650 ;
        RECT  7.410 0.470 8.810 0.590 ;
        RECT  7.290 0.470 7.410 0.830 ;
        RECT  6.580 0.710 7.290 0.830 ;
        RECT  6.580 1.450 6.740 1.610 ;
        RECT  6.460 0.710 6.580 1.610 ;
        RECT  10.660 1.050 10.890 1.270 ;
        RECT  10.540 1.050 10.660 2.050 ;
        RECT  9.130 1.930 10.540 2.050 ;
        RECT  9.010 1.770 9.130 2.050 ;
        RECT  8.490 1.770 9.010 1.890 ;
        RECT  8.490 1.050 8.520 1.270 ;
        RECT  8.370 0.710 8.490 1.890 ;
        RECT  7.530 0.710 8.370 0.870 ;
        RECT  6.230 0.810 6.460 0.970 ;
        RECT  7.140 1.620 8.370 1.780 ;
        RECT  5.900 0.760 6.060 1.280 ;
        RECT  3.690 1.930 3.930 2.090 ;
        RECT  4.090 1.300 4.330 1.460 ;
        RECT  3.860 0.430 4.030 0.590 ;
        RECT  3.510 1.650 3.630 1.810 ;
        RECT  3.890 1.650 4.420 1.810 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.850 1.500 3.050 1.660 ;
        RECT  2.160 1.640 2.610 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
        LAYER M1 ;
        RECT  10.830 1.650 10.935 2.030 ;
        RECT  10.830 0.490 10.935 0.870 ;
        RECT  9.450 0.490 9.655 0.870 ;
        RECT  9.430 1.600 9.655 1.760 ;
    END
END SDFNCSND4

MACRO SDFND1
    CLASS CORE ;
    FOREIGN SDFND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.720 1.960 7.750 2.100 ;
        RECT  7.750 0.420 7.910 2.100 ;
        RECT  7.910 1.960 7.940 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.890 1.960 6.920 2.100 ;
        RECT  6.920 1.390 7.080 2.100 ;
        RECT  7.080 1.960 7.110 2.100 ;
        RECT  7.080 1.390 7.130 1.515 ;
        RECT  6.920 0.710 7.130 0.870 ;
        RECT  7.130 0.710 7.270 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 2.710 0.300 ;
        RECT  2.710 -0.300 2.930 0.340 ;
        RECT  2.930 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.740 ;
        RECT  4.690 -0.300 6.150 0.300 ;
        RECT  6.150 -0.300 6.370 0.340 ;
        RECT  6.370 -0.300 7.320 0.300 ;
        RECT  7.320 -0.300 7.540 0.340 ;
        RECT  7.540 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.700 2.820 ;
        RECT  2.700 2.180 2.920 2.820 ;
        RECT  2.920 2.220 4.380 2.820 ;
        RECT  4.380 2.000 4.600 2.820 ;
        RECT  4.600 2.220 6.140 2.820 ;
        RECT  6.140 2.180 6.360 2.820 ;
        RECT  6.360 2.220 7.310 2.820 ;
        RECT  7.310 2.180 7.530 2.820 ;
        RECT  7.530 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.260 0.710 5.350 2.050 ;
        RECT  5.350 0.710 5.420 0.930 ;
        RECT  5.350 1.930 6.190 2.050 ;
        RECT  6.190 1.390 6.310 2.050 ;
        RECT  6.310 1.390 6.340 1.510 ;
        RECT  6.340 1.050 6.460 1.510 ;
        RECT  6.460 1.050 6.560 1.270 ;
        RECT  5.470 1.150 5.540 1.750 ;
        RECT  5.320 0.470 5.540 0.590 ;
        RECT  5.540 0.470 5.630 1.750 ;
        RECT  5.630 0.470 5.660 1.270 ;
        RECT  4.500 0.860 4.880 0.980 ;
        RECT  4.760 1.630 4.940 1.790 ;
        RECT  4.880 0.700 4.940 0.980 ;
        RECT  4.940 0.700 5.040 1.790 ;
        RECT  5.040 0.860 5.060 1.790 ;
        RECT  4.010 1.390 4.660 1.510 ;
        RECT  4.660 1.100 4.820 1.510 ;
        RECT  1.350 0.470 3.440 0.590 ;
        RECT  3.440 0.470 3.660 0.775 ;
        RECT  1.410 1.930 3.470 2.050 ;
        RECT  3.470 1.530 3.630 2.050 ;
        RECT  3.150 0.710 3.170 0.930 ;
        RECT  3.170 0.710 3.290 1.810 ;
        RECT  3.290 1.080 3.565 1.240 ;
        RECT  2.280 0.710 2.910 0.870 ;
        RECT  2.910 0.710 3.030 1.810 ;
        RECT  3.030 1.050 3.050 1.270 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.430 1.810 1.670 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  6.800 1.080 7.010 1.240 ;
        RECT  6.740 0.710 6.800 1.510 ;
        RECT  6.740 1.960 6.770 2.100 ;
        RECT  6.680 0.710 6.740 2.100 ;
        RECT  6.200 0.710 6.680 0.870 ;
        RECT  6.580 1.390 6.680 2.100 ;
        RECT  6.550 1.960 6.580 2.100 ;
        RECT  7.470 0.470 7.630 1.290 ;
        RECT  5.920 0.470 7.470 0.590 ;
        RECT  5.910 0.470 5.920 1.580 ;
        RECT  5.780 0.470 5.910 1.810 ;
        RECT  5.750 1.460 5.780 1.810 ;
        RECT  6.040 0.710 6.200 1.270 ;
        RECT  5.190 0.810 5.260 2.050 ;
        RECT  5.100 0.420 5.320 0.590 ;
        RECT  4.340 0.860 4.500 1.270 ;
        RECT  3.850 0.565 4.010 2.040 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.150 1.590 3.170 1.810 ;
        RECT  2.350 1.650 2.910 1.810 ;
        RECT  1.530 0.710 1.650 1.575 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFND1

MACRO SDFND2
    CLASS CORE ;
    FOREIGN SDFND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.000 1.960 8.030 2.100 ;
        RECT  8.030 1.390 8.090 2.100 ;
        RECT  8.030 0.420 8.090 0.900 ;
        RECT  8.090 0.420 8.190 2.100 ;
        RECT  8.190 1.960 8.220 2.100 ;
        RECT  8.190 0.780 8.230 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.220 1.960 7.250 2.100 ;
        RECT  7.250 1.390 7.410 2.100 ;
        RECT  7.410 1.960 7.440 2.100 ;
        RECT  7.410 1.390 7.450 1.515 ;
        RECT  7.230 0.710 7.450 0.870 ;
        RECT  7.450 0.710 7.590 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.950 0.300 ;
        RECT  1.950 -0.300 2.170 0.340 ;
        RECT  2.170 -0.300 2.680 0.300 ;
        RECT  2.680 -0.300 2.900 0.340 ;
        RECT  2.900 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.740 ;
        RECT  4.670 -0.300 6.130 0.300 ;
        RECT  6.130 -0.300 6.350 0.340 ;
        RECT  6.350 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.680 2.820 ;
        RECT  2.680 2.180 2.900 2.820 ;
        RECT  2.900 2.220 4.360 2.820 ;
        RECT  4.360 2.000 4.580 2.820 ;
        RECT  4.580 2.220 6.120 2.820 ;
        RECT  6.120 2.180 6.340 2.820 ;
        RECT  6.340 2.220 7.610 2.820 ;
        RECT  7.610 2.180 7.830 2.820 ;
        RECT  7.830 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.350 0.470 3.420 0.590 ;
        RECT  3.420 0.470 3.640 0.785 ;
        RECT  1.410 1.930 3.450 2.050 ;
        RECT  3.450 1.540 3.610 2.050 ;
        RECT  3.130 0.710 3.150 0.930 ;
        RECT  3.150 0.710 3.270 1.810 ;
        RECT  3.270 1.080 3.545 1.240 ;
        RECT  2.280 0.710 2.890 0.870 ;
        RECT  2.890 0.710 3.010 1.810 ;
        RECT  3.010 1.050 3.030 1.270 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.430 1.810 1.670 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  4.640 1.100 4.800 1.510 ;
        RECT  3.990 1.390 4.640 1.510 ;
        RECT  5.020 0.860 5.040 1.790 ;
        RECT  4.920 0.700 5.020 1.790 ;
        RECT  4.860 0.700 4.920 0.980 ;
        RECT  4.740 1.630 4.920 1.790 ;
        RECT  4.480 0.860 4.860 0.980 ;
        RECT  5.610 0.470 5.640 1.270 ;
        RECT  5.520 0.470 5.610 1.750 ;
        RECT  5.300 0.470 5.520 0.590 ;
        RECT  5.450 1.150 5.520 1.750 ;
        RECT  6.440 1.050 6.540 1.270 ;
        RECT  6.320 1.050 6.440 1.510 ;
        RECT  6.290 1.390 6.320 1.510 ;
        RECT  6.170 1.390 6.290 2.050 ;
        RECT  5.330 1.930 6.170 2.050 ;
        RECT  5.330 0.710 5.400 0.930 ;
        RECT  5.240 0.710 5.330 2.050 ;
        RECT  6.780 1.080 7.320 1.240 ;
        RECT  6.720 0.710 6.780 1.700 ;
        RECT  6.660 0.710 6.720 2.080 ;
        RECT  6.180 0.710 6.660 0.870 ;
        RECT  6.560 1.580 6.660 2.080 ;
        RECT  7.750 0.470 7.910 1.290 ;
        RECT  5.900 0.470 7.750 0.590 ;
        RECT  5.890 0.470 5.900 1.580 ;
        RECT  5.760 0.470 5.890 1.810 ;
        RECT  5.730 1.460 5.760 1.810 ;
        RECT  6.020 0.710 6.180 1.270 ;
        RECT  5.170 0.810 5.240 2.050 ;
        RECT  5.080 0.420 5.300 0.590 ;
        RECT  4.320 0.860 4.480 1.270 ;
        RECT  3.830 0.575 3.990 2.050 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.130 1.590 3.150 1.810 ;
        RECT  2.350 1.650 2.890 1.810 ;
        RECT  1.530 0.710 1.650 1.575 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFND2

MACRO SDFND4
    CLASS CORE ;
    FOREIGN SDFND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.910 1.650 9.230 2.030 ;
        RECT  8.910 0.490 9.230 0.870 ;
        RECT  9.230 0.490 9.650 2.030 ;
        RECT  9.650 1.650 9.820 2.030 ;
        RECT  9.650 0.490 9.820 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.530 1.650 7.950 2.030 ;
        RECT  7.510 0.710 7.950 0.870 ;
        RECT  7.950 0.710 8.370 2.030 ;
        RECT  8.370 1.650 8.440 2.030 ;
        RECT  8.370 0.710 8.460 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.600 1.270 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 4.280 0.300 ;
        RECT  4.280 -0.300 4.500 0.740 ;
        RECT  4.500 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 4.320 2.820 ;
        RECT  4.320 2.030 4.540 2.820 ;
        RECT  4.540 2.220 5.750 2.820 ;
        RECT  5.750 2.180 5.970 2.820 ;
        RECT  5.970 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  1.650 1.430 1.810 1.670 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  2.840 1.050 2.920 1.270 ;
        RECT  2.720 0.710 2.840 1.810 ;
        RECT  2.170 0.710 2.720 0.870 ;
        RECT  3.160 1.080 3.435 1.240 ;
        RECT  3.040 0.710 3.160 1.810 ;
        RECT  2.970 0.710 3.040 0.930 ;
        RECT  3.290 0.470 3.450 0.850 ;
        RECT  1.350 0.470 3.290 0.590 ;
        RECT  3.330 1.540 3.490 2.050 ;
        RECT  1.410 1.930 3.330 2.050 ;
        RECT  4.530 1.100 4.690 1.510 ;
        RECT  3.870 1.390 4.530 1.510 ;
        RECT  3.860 1.390 3.870 2.050 ;
        RECT  3.710 0.580 3.860 2.050 ;
        RECT  4.850 0.860 4.970 1.790 ;
        RECT  4.690 0.650 4.850 0.980 ;
        RECT  4.700 1.630 4.850 1.790 ;
        RECT  4.370 0.860 4.690 0.980 ;
        RECT  6.840 1.030 7.000 1.510 ;
        RECT  6.705 1.390 6.840 1.510 ;
        RECT  6.585 1.390 6.705 2.050 ;
        RECT  5.290 1.930 6.585 2.050 ;
        RECT  5.230 1.395 5.290 2.050 ;
        RECT  5.130 0.650 5.230 2.050 ;
        RECT  7.340 1.080 7.635 1.240 ;
        RECT  7.220 0.710 7.340 1.775 ;
        RECT  6.620 0.710 7.220 0.870 ;
        RECT  7.060 1.650 7.220 1.775 ;
        RECT  6.840 1.650 7.060 2.070 ;
        RECT  6.500 0.710 6.620 1.240 ;
        RECT  8.770 1.080 9.015 1.240 ;
        RECT  8.610 0.470 8.770 1.240 ;
        RECT  6.370 0.470 8.610 0.590 ;
        RECT  5.730 1.620 6.390 1.780 ;
        RECT  6.150 0.470 6.370 0.680 ;
        RECT  5.730 0.560 6.150 0.680 ;
        RECT  5.610 0.560 5.730 1.780 ;
        RECT  5.420 0.700 5.610 0.860 ;
        RECT  5.490 1.620 5.610 1.780 ;
        RECT  6.280 1.080 6.500 1.240 ;
        RECT  5.090 0.650 5.130 1.515 ;
        RECT  4.210 0.860 4.370 1.270 ;
        RECT  3.620 0.580 3.710 0.740 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  2.990 1.590 3.040 1.810 ;
        RECT  2.240 1.650 2.720 1.810 ;
        RECT  1.530 0.710 1.650 1.575 ;
        RECT  0.100 0.590 0.260 0.880 ;
        LAYER M1 ;
        RECT  8.910 1.650 9.015 2.030 ;
        RECT  8.910 0.490 9.015 0.870 ;
        RECT  7.530 1.650 7.735 2.030 ;
        RECT  7.510 0.710 7.735 0.870 ;
    END
END SDFND4

MACRO SDFNSND1
    CLASS CORE ;
    FOREIGN SDFNSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.360 1.940 8.390 2.100 ;
        RECT  8.390 1.390 8.410 2.100 ;
        RECT  8.390 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.550 2.100 ;
        RECT  8.550 1.940 8.580 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.940 7.670 2.100 ;
        RECT  7.670 1.390 7.770 2.100 ;
        RECT  7.670 0.710 7.770 0.930 ;
        RECT  7.770 0.710 7.830 2.100 ;
        RECT  7.830 1.940 7.860 2.100 ;
        RECT  7.830 0.710 7.910 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.570 0.300 ;
        RECT  2.570 -0.300 2.790 0.340 ;
        RECT  2.790 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.900 0.710 7.430 0.850 ;
        RECT  7.430 0.710 7.490 2.100 ;
        RECT  7.490 1.940 7.520 2.100 ;
        RECT  7.490 0.710 7.550 1.515 ;
        RECT  7.550 1.050 7.650 1.270 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  7.050 1.050 7.170 1.900 ;
        RECT  7.170 1.050 7.310 1.270 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  3.800 0.720 3.920 1.780 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  2.960 0.710 3.110 0.870 ;
        RECT  3.110 0.710 3.230 1.660 ;
        RECT  3.230 1.110 3.680 1.270 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  1.280 1.920 3.320 2.040 ;
        RECT  3.320 1.800 3.480 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.080 2.990 1.240 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  7.330 1.390 7.430 2.100 ;
        RECT  7.300 1.940 7.330 2.100 ;
        RECT  8.260 1.050 8.290 1.290 ;
        RECT  8.140 0.470 8.260 1.290 ;
        RECT  6.570 0.470 8.140 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.670 1.620 3.800 1.780 ;
        RECT  2.910 1.500 3.110 1.660 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  5.950 1.410 6.450 1.570 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFNSND1

MACRO SDFNSND2
    CLASS CORE ;
    FOREIGN SDFNSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.940 8.990 2.100 ;
        RECT  8.990 1.390 9.050 2.100 ;
        RECT  8.990 0.420 9.050 0.900 ;
        RECT  9.050 0.420 9.150 2.100 ;
        RECT  9.150 1.940 9.180 2.100 ;
        RECT  9.150 0.780 9.190 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.160 1.940 8.190 2.100 ;
        RECT  8.190 1.390 8.350 2.100 ;
        RECT  8.350 1.940 8.380 2.100 ;
        RECT  8.350 1.390 8.410 1.515 ;
        RECT  8.140 0.710 8.410 0.870 ;
        RECT  8.410 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.570 0.300 ;
        RECT  2.570 -0.300 2.790 0.340 ;
        RECT  2.790 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 7.760 0.300 ;
        RECT  7.760 -0.300 7.980 0.340 ;
        RECT  7.980 -0.300 8.560 0.300 ;
        RECT  8.560 -0.300 8.780 0.340 ;
        RECT  8.780 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.530 2.820 ;
        RECT  2.530 2.180 2.750 2.820 ;
        RECT  2.750 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 7.760 2.820 ;
        RECT  7.760 2.180 7.980 2.820 ;
        RECT  7.980 2.220 8.560 2.820 ;
        RECT  8.560 2.180 8.780 2.820 ;
        RECT  8.780 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  3.800 0.720 3.920 1.780 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  2.960 0.710 3.110 0.870 ;
        RECT  3.110 0.710 3.230 1.660 ;
        RECT  3.230 1.110 3.680 1.270 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  1.280 1.920 3.320 2.040 ;
        RECT  3.320 1.800 3.480 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.080 2.990 1.240 ;
        RECT  1.640 1.470 1.660 1.710 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  7.170 1.050 7.310 1.270 ;
        RECT  7.050 1.050 7.170 1.900 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  7.550 1.080 8.270 1.240 ;
        RECT  7.490 0.710 7.550 1.705 ;
        RECT  7.430 0.710 7.490 2.080 ;
        RECT  6.900 0.710 7.430 0.850 ;
        RECT  7.330 1.580 7.430 2.080 ;
        RECT  8.870 1.050 8.930 1.270 ;
        RECT  8.750 0.470 8.870 1.270 ;
        RECT  6.570 0.470 8.750 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  5.950 1.410 6.450 1.570 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.670 1.620 3.800 1.780 ;
        RECT  2.910 1.500 3.110 1.660 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.710 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFNSND2

MACRO SDFNSND4
    CLASS CORE ;
    FOREIGN SDFNSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.460 1.650 9.870 2.030 ;
        RECT  9.460 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 2.030 ;
        RECT  10.290 1.650 10.410 2.030 ;
        RECT  10.290 0.490 10.410 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.020 1.650 8.270 2.030 ;
        RECT  8.000 0.760 8.270 0.920 ;
        RECT  8.270 0.760 8.690 2.030 ;
        RECT  8.690 1.650 8.970 2.030 ;
        RECT  8.690 0.760 8.990 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CPN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.280 1.920 3.320 2.040 ;
        RECT  3.320 1.800 3.480 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.080 2.990 1.240 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  3.230 1.110 3.680 1.270 ;
        RECT  3.110 0.710 3.230 1.660 ;
        RECT  2.960 0.710 3.110 0.870 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  3.800 0.720 3.920 1.780 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  7.170 1.050 7.310 1.270 ;
        RECT  7.050 1.050 7.170 1.900 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  7.550 1.050 8.040 1.270 ;
        RECT  7.490 0.710 7.550 1.515 ;
        RECT  7.490 1.940 7.520 2.100 ;
        RECT  7.430 0.710 7.490 2.100 ;
        RECT  6.900 0.710 7.430 0.850 ;
        RECT  7.330 1.390 7.430 2.100 ;
        RECT  7.300 1.940 7.330 2.100 ;
        RECT  9.280 1.080 9.570 1.240 ;
        RECT  9.160 0.470 9.280 1.240 ;
        RECT  6.570 0.470 9.160 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  5.950 1.410 6.450 1.570 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.670 1.620 3.800 1.780 ;
        RECT  2.910 1.500 3.110 1.660 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
        LAYER M1 ;
        RECT  9.460 1.650 9.655 2.030 ;
        RECT  9.460 0.490 9.655 0.870 ;
        RECT  8.905 1.650 8.970 2.030 ;
        RECT  8.905 0.760 8.990 0.920 ;
        RECT  8.020 1.650 8.055 2.030 ;
        RECT  8.000 0.760 8.055 0.920 ;
    END
END SDFNSND4

MACRO SDFQD1
    CLASS CORE ;
    FOREIGN SDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.680 1.960 6.710 2.100 ;
        RECT  6.710 1.390 6.870 2.100 ;
        RECT  6.870 1.960 6.900 2.100 ;
        RECT  6.710 0.450 6.930 0.870 ;
        RECT  6.870 1.390 7.130 1.515 ;
        RECT  6.930 0.710 7.130 0.870 ;
        RECT  7.130 0.710 7.270 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.700 0.300 ;
        RECT  2.700 -0.300 2.920 0.340 ;
        RECT  2.920 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.740 ;
        RECT  4.690 -0.300 5.950 0.300 ;
        RECT  5.950 -0.300 6.170 0.340 ;
        RECT  6.170 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.700 2.820 ;
        RECT  2.700 2.180 2.920 2.820 ;
        RECT  2.920 2.220 4.480 2.820 ;
        RECT  4.480 2.000 4.700 2.820 ;
        RECT  4.700 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.660 1.340 5.730 1.750 ;
        RECT  4.500 0.860 4.880 0.980 ;
        RECT  4.860 1.630 4.980 1.790 ;
        RECT  4.880 0.700 4.980 0.980 ;
        RECT  4.980 0.700 5.040 1.790 ;
        RECT  5.040 0.860 5.100 1.790 ;
        RECT  4.010 1.390 4.680 1.510 ;
        RECT  4.680 1.100 4.840 1.510 ;
        RECT  1.350 0.470 3.440 0.590 ;
        RECT  3.440 0.470 3.680 0.630 ;
        RECT  1.410 1.930 3.470 2.050 ;
        RECT  3.470 1.420 3.630 2.050 ;
        RECT  3.150 0.710 3.170 0.930 ;
        RECT  3.170 0.710 3.290 1.810 ;
        RECT  3.290 1.080 3.565 1.240 ;
        RECT  2.270 0.710 2.910 0.870 ;
        RECT  2.910 0.710 3.030 1.810 ;
        RECT  3.030 1.050 3.050 1.270 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.460 1.860 1.620 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  5.570 0.470 5.660 1.750 ;
        RECT  5.540 0.470 5.570 1.460 ;
        RECT  5.320 0.470 5.540 0.590 ;
        RECT  6.250 1.050 6.350 1.270 ;
        RECT  6.130 1.050 6.250 1.510 ;
        RECT  6.100 1.390 6.130 1.510 ;
        RECT  5.980 1.390 6.100 2.050 ;
        RECT  5.450 1.930 5.980 2.050 ;
        RECT  5.420 1.570 5.450 2.050 ;
        RECT  5.290 0.710 5.420 2.050 ;
        RECT  6.590 1.080 7.010 1.240 ;
        RECT  6.570 0.710 6.590 1.510 ;
        RECT  6.530 0.450 6.570 1.510 ;
        RECT  6.530 1.960 6.560 2.100 ;
        RECT  6.470 0.450 6.530 2.100 ;
        RECT  6.350 0.450 6.470 0.870 ;
        RECT  6.370 1.390 6.470 2.100 ;
        RECT  6.340 1.960 6.370 2.100 ;
        RECT  5.990 0.710 6.350 0.870 ;
        RECT  5.830 0.710 5.990 1.270 ;
        RECT  5.260 0.710 5.290 1.690 ;
        RECT  5.100 0.420 5.320 0.590 ;
        RECT  4.340 0.860 4.500 1.270 ;
        RECT  3.850 0.450 4.010 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.150 1.590 3.170 1.810 ;
        RECT  2.350 1.650 2.910 1.810 ;
        RECT  1.530 0.710 1.650 1.620 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFQD1

MACRO SDFQD2
    CLASS CORE ;
    FOREIGN SDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.030 1.960 7.060 2.100 ;
        RECT  7.060 1.390 7.220 2.100 ;
        RECT  7.060 0.420 7.220 0.900 ;
        RECT  7.220 1.960 7.250 2.100 ;
        RECT  7.220 1.390 7.450 1.515 ;
        RECT  7.220 0.770 7.450 0.900 ;
        RECT  7.450 0.770 7.590 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.730 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.930 0.300 ;
        RECT  1.930 -0.300 2.150 0.340 ;
        RECT  2.150 -0.300 2.700 0.300 ;
        RECT  2.700 -0.300 2.920 0.340 ;
        RECT  2.920 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.740 ;
        RECT  4.690 -0.300 5.940 0.300 ;
        RECT  5.940 -0.300 6.160 0.340 ;
        RECT  6.160 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 2.020 2.820 ;
        RECT  2.020 2.180 2.240 2.820 ;
        RECT  2.240 2.220 2.700 2.820 ;
        RECT  2.700 2.180 2.920 2.820 ;
        RECT  2.920 2.220 4.480 2.820 ;
        RECT  4.480 2.000 4.700 2.820 ;
        RECT  4.700 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  1.650 1.460 1.860 1.620 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  3.030 1.050 3.050 1.270 ;
        RECT  2.910 0.710 3.030 1.810 ;
        RECT  2.270 0.710 2.910 0.870 ;
        RECT  3.290 1.080 3.565 1.240 ;
        RECT  3.170 0.710 3.290 1.810 ;
        RECT  3.150 0.710 3.170 0.930 ;
        RECT  3.470 1.420 3.630 2.050 ;
        RECT  1.410 1.930 3.470 2.050 ;
        RECT  3.440 0.470 3.680 0.630 ;
        RECT  1.350 0.470 3.440 0.590 ;
        RECT  4.680 1.100 4.840 1.510 ;
        RECT  4.010 1.390 4.680 1.510 ;
        RECT  5.040 0.860 5.100 1.790 ;
        RECT  4.980 0.700 5.040 1.790 ;
        RECT  4.880 0.700 4.980 0.980 ;
        RECT  4.860 1.630 4.980 1.790 ;
        RECT  4.500 0.860 4.880 0.980 ;
        RECT  5.660 1.340 5.730 1.750 ;
        RECT  5.570 0.470 5.660 1.750 ;
        RECT  5.540 0.470 5.570 1.460 ;
        RECT  5.320 0.470 5.540 0.590 ;
        RECT  6.250 1.050 6.350 1.270 ;
        RECT  6.130 1.050 6.250 1.510 ;
        RECT  6.100 1.390 6.130 1.510 ;
        RECT  5.980 1.390 6.100 2.050 ;
        RECT  5.450 1.930 5.980 2.050 ;
        RECT  5.420 1.570 5.450 2.050 ;
        RECT  5.290 0.710 5.420 2.050 ;
        RECT  6.590 1.080 7.190 1.240 ;
        RECT  6.530 0.710 6.590 1.700 ;
        RECT  6.470 0.710 6.530 2.080 ;
        RECT  5.990 0.710 6.470 0.870 ;
        RECT  6.370 1.580 6.470 2.080 ;
        RECT  5.260 0.710 5.290 1.690 ;
        RECT  5.100 0.420 5.320 0.590 ;
        RECT  4.340 0.860 4.500 1.270 ;
        RECT  3.850 0.450 4.010 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.150 1.590 3.170 1.810 ;
        RECT  2.350 1.650 2.910 1.810 ;
        RECT  1.530 0.710 1.650 1.620 ;
        RECT  5.830 0.710 5.990 1.270 ;
        RECT  0.100 0.590 0.260 0.880 ;
    END
END SDFQD2

MACRO SDFQD4
    CLASS CORE ;
    FOREIGN SDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.990 1.650 7.310 2.030 ;
        RECT  6.990 0.490 7.310 0.870 ;
        RECT  7.310 0.490 7.730 2.030 ;
        RECT  7.730 1.650 7.900 2.030 ;
        RECT  7.730 0.490 7.900 0.870 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.790 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.005 2.470 1.515 ;
        RECT  2.470 1.050 2.690 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.470 0.300 ;
        RECT  0.470 -0.300 0.690 0.640 ;
        RECT  0.690 -0.300 1.920 0.300 ;
        RECT  1.920 -0.300 2.140 0.340 ;
        RECT  2.140 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.890 0.340 ;
        RECT  2.890 -0.300 4.430 0.300 ;
        RECT  4.430 -0.300 4.650 0.740 ;
        RECT  4.650 -0.300 5.900 0.300 ;
        RECT  5.900 -0.300 6.120 0.340 ;
        RECT  6.120 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.950 0.690 2.820 ;
        RECT  0.690 2.220 4.440 2.820 ;
        RECT  4.440 2.000 4.660 2.820 ;
        RECT  4.660 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.830 ;
        RECT  0.490 0.760 1.090 0.880 ;
        RECT  1.090 0.760 1.250 1.420 ;
        RECT  0.070 1.670 0.370 1.830 ;
        RECT  1.650 1.460 1.860 1.620 ;
        RECT  1.650 0.710 1.770 0.870 ;
        RECT  2.990 1.050 3.010 1.270 ;
        RECT  2.870 0.710 2.990 1.810 ;
        RECT  2.240 0.710 2.870 0.870 ;
        RECT  3.250 1.080 3.525 1.240 ;
        RECT  3.130 0.710 3.250 1.810 ;
        RECT  3.110 0.710 3.130 0.930 ;
        RECT  3.430 1.420 3.590 2.050 ;
        RECT  1.410 1.930 3.430 2.050 ;
        RECT  3.400 0.470 3.640 0.630 ;
        RECT  1.350 0.470 3.400 0.590 ;
        RECT  4.640 1.100 4.800 1.510 ;
        RECT  3.970 1.390 4.640 1.510 ;
        RECT  5.000 0.860 5.060 1.790 ;
        RECT  4.940 0.700 5.000 1.790 ;
        RECT  4.840 0.700 4.940 0.980 ;
        RECT  4.820 1.630 4.940 1.790 ;
        RECT  4.460 0.860 4.840 0.980 ;
        RECT  5.620 1.340 5.690 1.750 ;
        RECT  5.530 0.470 5.620 1.750 ;
        RECT  5.500 0.470 5.530 1.460 ;
        RECT  5.280 0.470 5.500 0.590 ;
        RECT  6.210 1.080 6.370 1.240 ;
        RECT  6.090 1.080 6.210 1.510 ;
        RECT  6.060 1.390 6.090 1.510 ;
        RECT  5.940 1.390 6.060 2.050 ;
        RECT  5.410 1.930 5.940 2.050 ;
        RECT  5.380 1.570 5.410 2.050 ;
        RECT  5.250 0.710 5.380 2.050 ;
        RECT  6.610 1.080 7.095 1.240 ;
        RECT  6.490 0.760 6.610 1.500 ;
        RECT  6.490 1.930 6.520 2.090 ;
        RECT  6.330 0.420 6.490 0.920 ;
        RECT  6.330 1.380 6.490 2.090 ;
        RECT  5.950 0.760 6.330 0.920 ;
        RECT  6.300 1.930 6.330 2.090 ;
        RECT  5.220 0.710 5.250 1.690 ;
        RECT  5.060 0.420 5.280 0.590 ;
        RECT  4.300 0.860 4.460 1.270 ;
        RECT  3.810 0.450 3.970 1.930 ;
        RECT  1.110 0.470 1.350 0.630 ;
        RECT  1.250 1.620 1.410 2.050 ;
        RECT  3.110 1.590 3.130 1.810 ;
        RECT  2.310 1.650 2.870 1.810 ;
        RECT  1.530 0.710 1.650 1.620 ;
        RECT  5.790 0.760 5.950 1.270 ;
        RECT  0.100 0.590 0.260 0.880 ;
        LAYER M1 ;
        RECT  6.990 1.650 7.095 2.030 ;
        RECT  6.990 0.490 7.095 0.870 ;
    END
END SDFQD4

MACRO SDFSND1
    CLASS CORE ;
    FOREIGN SDFSND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.360 1.940 8.390 2.100 ;
        RECT  8.390 1.390 8.410 2.100 ;
        RECT  8.390 0.420 8.410 0.900 ;
        RECT  8.410 0.420 8.550 2.100 ;
        RECT  8.550 1.940 8.580 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  7.640 1.940 7.670 2.100 ;
        RECT  7.670 1.390 7.770 2.100 ;
        RECT  7.670 0.710 7.770 0.930 ;
        RECT  7.770 0.710 7.830 2.100 ;
        RECT  7.830 1.940 7.860 2.100 ;
        RECT  7.830 0.710 7.910 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.570 0.300 ;
        RECT  2.570 -0.300 2.790 0.340 ;
        RECT  2.790 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 8.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 8.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.900 0.710 7.430 0.850 ;
        RECT  7.430 0.710 7.490 2.100 ;
        RECT  7.490 1.940 7.520 2.100 ;
        RECT  7.490 0.710 7.550 1.515 ;
        RECT  7.550 1.050 7.650 1.270 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  7.050 1.050 7.170 1.900 ;
        RECT  7.170 1.050 7.310 1.270 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  3.800 0.720 3.920 1.750 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  2.960 0.710 3.090 0.870 ;
        RECT  3.090 0.710 3.210 1.660 ;
        RECT  3.210 1.110 3.460 1.270 ;
        RECT  1.280 1.920 3.300 2.040 ;
        RECT  3.300 1.745 3.460 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.050 2.960 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  7.330 1.390 7.430 2.100 ;
        RECT  7.300 1.940 7.330 2.100 ;
        RECT  8.260 1.050 8.290 1.290 ;
        RECT  8.140 0.470 8.260 1.290 ;
        RECT  6.570 0.470 8.140 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.650 1.590 3.800 1.750 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.890 1.500 3.090 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
        RECT  5.950 1.410 6.450 1.570 ;
    END
END SDFSND1

MACRO SDFSND2
    CLASS CORE ;
    FOREIGN SDFSND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.940 8.990 2.100 ;
        RECT  8.990 1.390 9.050 2.100 ;
        RECT  8.990 0.420 9.050 0.900 ;
        RECT  9.050 0.420 9.150 2.100 ;
        RECT  9.150 1.940 9.180 2.100 ;
        RECT  9.150 0.780 9.190 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.260 1.940 8.290 2.100 ;
        RECT  8.290 1.390 8.410 2.100 ;
        RECT  8.240 0.710 8.410 0.870 ;
        RECT  8.410 0.710 8.450 2.100 ;
        RECT  8.450 1.940 8.480 2.100 ;
        RECT  8.450 0.710 8.550 1.515 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 1.980 0.300 ;
        RECT  1.980 -0.300 2.200 0.340 ;
        RECT  2.200 -0.300 2.570 0.300 ;
        RECT  2.570 -0.300 2.790 0.340 ;
        RECT  2.790 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 7.860 0.300 ;
        RECT  7.860 -0.300 8.080 0.340 ;
        RECT  8.080 -0.300 9.600 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 2.510 2.820 ;
        RECT  2.510 2.180 2.730 2.820 ;
        RECT  2.730 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 7.010 2.820 ;
        RECT  7.010 2.180 7.230 2.820 ;
        RECT  7.230 2.220 7.860 2.820 ;
        RECT  7.860 2.180 8.080 2.820 ;
        RECT  8.080 2.220 9.600 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.960 0.710 3.090 0.870 ;
        RECT  3.090 0.710 3.210 1.660 ;
        RECT  3.210 1.110 3.460 1.270 ;
        RECT  1.280 1.920 3.300 2.040 ;
        RECT  3.300 1.745 3.460 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.050 2.960 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  3.800 0.720 3.920 1.750 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  7.170 1.080 7.420 1.240 ;
        RECT  7.050 1.080 7.170 1.900 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  7.660 1.050 8.260 1.270 ;
        RECT  7.600 0.710 7.660 1.745 ;
        RECT  7.540 0.710 7.600 2.100 ;
        RECT  6.900 0.710 7.540 0.850 ;
        RECT  7.440 1.620 7.540 2.100 ;
        RECT  8.845 1.050 8.930 1.270 ;
        RECT  8.725 0.470 8.845 1.270 ;
        RECT  6.570 0.470 8.725 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.650 1.590 3.800 1.750 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.890 1.500 3.090 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  5.950 1.410 6.450 1.570 ;
        RECT  0.080 0.760 0.100 1.850 ;
    END
END SDFSND2

MACRO SDFSND4
    CLASS CORE ;
    FOREIGN SDFSND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.670 1.050 0.730 1.270 ;
        RECT  0.730 1.005 0.870 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.330 1.050 0.410 1.270 ;
        RECT  0.410 1.005 0.550 1.515 ;
        END
    END SE
    PIN SDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.040 1.230 5.210 1.390 ;
        RECT  5.210 0.725 5.350 1.390 ;
        END
    END SDN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.460 1.650 9.870 2.030 ;
        RECT  9.460 0.490 9.870 0.870 ;
        RECT  9.870 0.490 10.290 2.030 ;
        RECT  10.290 1.650 10.410 2.030 ;
        RECT  10.290 0.490 10.410 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  8.020 1.650 8.270 2.030 ;
        RECT  8.000 0.760 8.270 0.920 ;
        RECT  8.270 0.760 8.690 2.030 ;
        RECT  8.690 1.650 8.970 2.030 ;
        RECT  8.690 0.760 8.990 0.920 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.775 1.050 2.010 1.270 ;
        RECT  2.010 1.005 2.150 1.515 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.460 0.300 ;
        RECT  0.460 -0.300 0.680 0.640 ;
        RECT  0.680 -0.300 4.270 0.300 ;
        RECT  4.270 -0.300 4.490 0.340 ;
        RECT  4.490 -0.300 6.890 0.300 ;
        RECT  6.890 -0.300 7.110 0.340 ;
        RECT  7.110 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.640 0.680 2.820 ;
        RECT  0.680 2.220 1.870 2.820 ;
        RECT  1.870 2.180 2.090 2.820 ;
        RECT  2.090 2.220 4.230 2.820 ;
        RECT  4.230 2.180 4.450 2.820 ;
        RECT  4.450 2.220 5.040 2.820 ;
        RECT  5.040 2.050 5.260 2.820 ;
        RECT  5.260 2.220 6.210 2.820 ;
        RECT  6.210 2.020 6.430 2.820 ;
        RECT  6.430 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.280 1.920 3.300 2.040 ;
        RECT  3.300 1.745 3.460 2.040 ;
        RECT  2.270 0.710 2.650 0.870 ;
        RECT  2.650 0.710 2.770 1.800 ;
        RECT  2.770 1.050 2.960 1.270 ;
        RECT  1.640 1.480 1.660 1.720 ;
        RECT  1.640 0.710 1.800 0.870 ;
        RECT  0.100 0.590 0.200 1.850 ;
        RECT  0.200 0.590 0.260 0.880 ;
        RECT  0.200 1.690 0.320 1.850 ;
        RECT  0.260 0.760 0.990 0.880 ;
        RECT  0.990 0.760 1.130 1.290 ;
        RECT  3.210 1.110 3.460 1.270 ;
        RECT  3.090 0.710 3.210 1.660 ;
        RECT  2.960 0.710 3.090 0.870 ;
        RECT  3.350 0.470 3.510 0.880 ;
        RECT  1.380 0.470 3.350 0.590 ;
        RECT  4.520 1.190 4.680 1.430 ;
        RECT  3.920 1.310 4.520 1.430 ;
        RECT  3.800 0.720 3.920 1.750 ;
        RECT  3.680 0.720 3.800 0.880 ;
        RECT  4.920 1.550 5.520 1.690 ;
        RECT  4.950 0.710 5.090 0.930 ;
        RECT  4.920 0.810 4.950 0.930 ;
        RECT  4.800 0.810 4.920 1.690 ;
        RECT  4.360 0.810 4.800 0.930 ;
        RECT  4.620 1.550 4.800 1.690 ;
        RECT  5.425 1.810 5.585 2.100 ;
        RECT  4.160 1.810 5.425 1.930 ;
        RECT  4.040 1.810 4.160 2.070 ;
        RECT  5.960 0.430 6.200 0.590 ;
        RECT  4.100 0.470 5.960 0.590 ;
        RECT  7.170 1.050 7.270 1.270 ;
        RECT  7.050 1.050 7.170 1.900 ;
        RECT  5.870 1.780 7.050 1.900 ;
        RECT  5.830 1.780 5.870 2.070 ;
        RECT  5.710 1.310 5.830 2.070 ;
        RECT  5.610 1.310 5.710 1.430 ;
        RECT  7.550 1.050 8.040 1.270 ;
        RECT  7.490 0.710 7.550 1.515 ;
        RECT  7.490 1.940 7.520 2.100 ;
        RECT  7.430 0.710 7.490 2.100 ;
        RECT  6.900 0.710 7.430 0.850 ;
        RECT  7.330 1.390 7.430 2.100 ;
        RECT  7.300 1.940 7.330 2.100 ;
        RECT  9.265 1.080 9.570 1.240 ;
        RECT  9.145 0.470 9.265 1.240 ;
        RECT  6.570 0.470 9.145 0.590 ;
        RECT  6.570 1.500 6.850 1.660 ;
        RECT  6.450 0.470 6.570 1.660 ;
        RECT  5.780 0.740 6.450 0.900 ;
        RECT  6.740 0.710 6.900 1.290 ;
        RECT  5.470 0.710 5.610 1.430 ;
        RECT  3.860 0.430 4.100 0.590 ;
        RECT  3.830 1.910 4.040 2.070 ;
        RECT  4.200 0.810 4.360 1.190 ;
        RECT  3.650 1.590 3.800 1.750 ;
        RECT  1.140 0.430 1.380 0.590 ;
        RECT  2.890 1.500 3.090 1.660 ;
        RECT  1.120 1.580 1.280 2.040 ;
        RECT  2.200 1.640 2.650 1.800 ;
        RECT  1.500 0.710 1.640 1.720 ;
        RECT  0.080 0.760 0.100 1.850 ;
        RECT  5.950 1.410 6.450 1.570 ;
        LAYER M1 ;
        RECT  9.460 1.650 9.655 2.030 ;
        RECT  9.460 0.490 9.655 0.870 ;
        RECT  8.905 1.650 8.970 2.030 ;
        RECT  8.905 0.760 8.990 0.920 ;
        RECT  8.020 1.650 8.055 2.030 ;
        RECT  8.000 0.760 8.055 0.920 ;
    END
END SDFSND4

MACRO SDFXD1
    CLASS CORE ;
    FOREIGN SDFXD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.240 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.270 3.110 1.795 ;
        RECT  3.110 1.270 3.150 1.510 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.380 3.930 1.540 ;
        RECT  3.930 1.005 4.070 1.540 ;
        END
    END SE
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.980 1.570 10.010 2.070 ;
        RECT  9.980 0.420 10.010 0.920 ;
        RECT  10.010 0.420 10.140 2.070 ;
        RECT  10.140 0.800 10.150 1.690 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.130 1.650 9.370 1.810 ;
        RECT  9.130 0.740 9.370 0.900 ;
        RECT  9.370 0.740 9.510 1.810 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.110 1.370 1.330 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 4.710 1.515 ;
        RECT  4.710 1.050 4.900 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 2.800 0.300 ;
        RECT  2.800 -0.300 3.020 0.760 ;
        RECT  3.020 -0.300 4.250 0.300 ;
        RECT  4.250 -0.300 4.470 0.340 ;
        RECT  4.470 -0.300 4.850 0.300 ;
        RECT  4.850 -0.300 5.070 0.340 ;
        RECT  5.070 -0.300 6.540 0.300 ;
        RECT  6.540 -0.300 6.760 0.760 ;
        RECT  6.760 -0.300 9.550 0.300 ;
        RECT  9.550 -0.300 9.770 0.340 ;
        RECT  9.770 -0.300 10.240 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.800 2.820 ;
        RECT  2.800 1.920 3.020 2.820 ;
        RECT  3.020 2.220 4.370 2.820 ;
        RECT  4.370 2.180 4.590 2.820 ;
        RECT  4.590 2.220 4.910 2.820 ;
        RECT  4.910 2.180 5.130 2.820 ;
        RECT  5.130 2.220 6.520 2.820 ;
        RECT  6.520 2.030 6.740 2.820 ;
        RECT  6.740 2.220 8.190 2.820 ;
        RECT  8.190 2.180 8.410 2.820 ;
        RECT  8.410 2.220 9.550 2.820 ;
        RECT  9.550 2.180 9.770 2.820 ;
        RECT  9.770 2.220 10.240 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.640 0.470 5.520 0.590 ;
        RECT  5.520 0.420 5.760 0.590 ;
        RECT  4.500 0.710 5.030 0.870 ;
        RECT  5.030 0.710 5.150 1.800 ;
        RECT  5.150 1.050 5.280 1.270 ;
        RECT  3.830 0.710 4.190 0.870 ;
        RECT  4.190 0.710 4.310 1.800 ;
        RECT  2.600 0.910 3.460 1.070 ;
        RECT  3.460 0.910 3.620 1.560 ;
        RECT  2.110 0.470 2.160 0.690 ;
        RECT  2.160 0.470 2.280 1.780 ;
        RECT  2.280 0.470 2.560 0.630 ;
        RECT  1.820 1.190 1.870 1.800 ;
        RECT  1.070 0.470 1.870 0.630 ;
        RECT  1.870 0.470 1.940 1.800 ;
        RECT  1.940 0.470 1.990 1.350 ;
        RECT  1.990 1.190 2.040 1.350 ;
        RECT  0.060 0.470 0.650 0.630 ;
        RECT  0.650 0.470 0.810 1.800 ;
        RECT  0.810 0.750 1.630 0.870 ;
        RECT  1.630 0.750 1.750 1.050 ;
        RECT  5.580 1.920 5.820 2.080 ;
        RECT  3.760 1.920 5.580 2.040 ;
        RECT  5.520 1.120 6.040 1.280 ;
        RECT  5.400 0.710 5.520 1.760 ;
        RECT  5.300 0.710 5.400 0.930 ;
        RECT  6.830 1.170 6.880 1.410 ;
        RECT  6.710 1.170 6.830 1.690 ;
        RECT  6.280 1.570 6.710 1.690 ;
        RECT  6.160 0.610 6.280 1.690 ;
        RECT  5.890 0.610 6.160 0.770 ;
        RECT  7.000 0.530 7.120 1.930 ;
        RECT  6.950 0.530 7.000 1.040 ;
        RECT  6.950 1.690 7.000 1.930 ;
        RECT  8.590 1.050 8.750 1.480 ;
        RECT  7.490 1.360 8.590 1.480 ;
        RECT  8.990 1.050 9.250 1.270 ;
        RECT  8.870 0.710 8.990 1.810 ;
        RECT  8.820 0.710 8.870 0.930 ;
        RECT  8.740 1.650 8.870 1.810 ;
        RECT  8.440 0.810 8.820 0.930 ;
        RECT  8.320 0.810 8.440 1.240 ;
        RECT  9.770 1.050 9.890 1.270 ;
        RECT  9.650 0.470 9.770 2.050 ;
        RECT  8.310 0.470 9.650 0.590 ;
        RECT  8.450 1.930 9.650 2.050 ;
        RECT  8.330 1.720 8.450 2.050 ;
        RECT  7.660 1.720 8.330 1.880 ;
        RECT  7.870 0.470 8.310 0.630 ;
        RECT  8.200 1.080 8.320 1.240 ;
        RECT  7.330 0.545 7.490 1.930 ;
        RECT  6.410 0.880 6.950 1.040 ;
        RECT  5.950 1.530 6.160 1.690 ;
        RECT  5.340 1.520 5.400 1.760 ;
        RECT  3.600 1.680 3.760 2.040 ;
        RECT  3.480 0.470 3.640 0.790 ;
        RECT  4.600 1.640 5.030 1.800 ;
        RECT  3.930 1.660 4.190 1.800 ;
        RECT  7.710 0.470 7.870 0.805 ;
        RECT  2.440 0.780 2.600 1.950 ;
        RECT  2.060 1.620 2.160 1.780 ;
        RECT  1.080 1.640 1.820 1.800 ;
        RECT  0.060 1.640 0.650 1.800 ;
    END
END SDFXD1

MACRO SDFXD2
    CLASS CORE ;
    FOREIGN SDFXD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.270 3.110 1.795 ;
        RECT  3.110 1.270 3.150 1.510 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.380 3.930 1.540 ;
        RECT  3.930 1.005 4.070 1.540 ;
        END
    END SE
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.210 1.570 10.370 2.070 ;
        RECT  10.210 0.420 10.370 0.920 ;
        RECT  10.370 1.570 10.650 1.690 ;
        RECT  10.370 0.800 10.650 0.920 ;
        RECT  10.650 0.800 10.790 1.690 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.430 1.635 9.690 1.795 ;
        RECT  9.450 0.760 9.690 0.920 ;
        RECT  9.690 0.760 9.830 1.795 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.110 1.370 1.330 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 4.710 1.515 ;
        RECT  4.710 1.050 4.900 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 2.800 0.300 ;
        RECT  2.800 -0.300 3.020 0.760 ;
        RECT  3.020 -0.300 4.250 0.300 ;
        RECT  4.250 -0.300 4.470 0.340 ;
        RECT  4.470 -0.300 4.850 0.300 ;
        RECT  4.850 -0.300 5.070 0.340 ;
        RECT  5.070 -0.300 6.540 0.300 ;
        RECT  6.540 -0.300 6.760 0.760 ;
        RECT  6.760 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.800 2.820 ;
        RECT  2.800 1.920 3.020 2.820 ;
        RECT  3.020 2.220 4.370 2.820 ;
        RECT  4.370 2.180 4.590 2.820 ;
        RECT  4.590 2.220 4.910 2.820 ;
        RECT  4.910 2.180 5.130 2.820 ;
        RECT  5.130 2.220 6.520 2.820 ;
        RECT  6.520 2.030 6.740 2.820 ;
        RECT  6.740 2.220 8.190 2.820 ;
        RECT  8.190 2.180 8.410 2.820 ;
        RECT  8.410 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.190 0.710 4.310 1.800 ;
        RECT  2.600 0.910 3.460 1.070 ;
        RECT  3.460 0.910 3.620 1.560 ;
        RECT  2.110 0.470 2.160 0.690 ;
        RECT  2.160 0.470 2.280 1.780 ;
        RECT  2.280 0.470 2.560 0.630 ;
        RECT  1.820 1.190 1.870 1.800 ;
        RECT  1.070 0.470 1.870 0.630 ;
        RECT  1.870 0.470 1.940 1.800 ;
        RECT  1.940 0.470 1.990 1.350 ;
        RECT  1.990 1.190 2.040 1.350 ;
        RECT  0.060 0.470 0.650 0.630 ;
        RECT  0.650 0.470 0.810 1.800 ;
        RECT  0.810 0.750 1.630 0.870 ;
        RECT  1.630 0.750 1.750 1.050 ;
        RECT  3.830 0.710 4.190 0.870 ;
        RECT  5.150 1.050 5.280 1.270 ;
        RECT  5.030 0.710 5.150 1.800 ;
        RECT  4.500 0.710 5.030 0.870 ;
        RECT  5.520 0.420 5.760 0.590 ;
        RECT  3.640 0.470 5.520 0.590 ;
        RECT  5.580 1.920 5.820 2.080 ;
        RECT  3.760 1.920 5.580 2.040 ;
        RECT  5.520 1.120 6.040 1.280 ;
        RECT  5.400 0.710 5.520 1.760 ;
        RECT  5.300 0.710 5.400 0.930 ;
        RECT  6.830 1.170 6.880 1.410 ;
        RECT  6.710 1.170 6.830 1.690 ;
        RECT  6.280 1.570 6.710 1.690 ;
        RECT  6.160 0.610 6.280 1.690 ;
        RECT  5.890 0.610 6.160 0.770 ;
        RECT  7.000 0.530 7.120 1.930 ;
        RECT  6.950 0.530 7.000 1.040 ;
        RECT  6.950 1.690 7.000 1.930 ;
        RECT  8.730 1.050 8.890 1.480 ;
        RECT  7.490 1.360 8.730 1.480 ;
        RECT  9.185 1.080 9.560 1.240 ;
        RECT  9.065 0.810 9.185 1.810 ;
        RECT  9.000 0.810 9.065 0.930 ;
        RECT  8.740 1.650 9.065 1.810 ;
        RECT  8.780 0.710 9.000 0.930 ;
        RECT  8.440 0.810 8.780 0.930 ;
        RECT  8.320 0.810 8.440 1.240 ;
        RECT  10.090 1.080 10.290 1.240 ;
        RECT  9.970 0.470 10.090 2.050 ;
        RECT  8.310 0.470 9.970 0.590 ;
        RECT  8.260 1.930 9.970 2.050 ;
        RECT  7.870 0.470 8.310 0.630 ;
        RECT  8.140 1.720 8.260 2.050 ;
        RECT  7.660 1.720 8.140 1.880 ;
        RECT  7.710 0.470 7.870 0.805 ;
        RECT  8.200 1.080 8.320 1.240 ;
        RECT  7.330 0.545 7.490 1.930 ;
        RECT  6.410 0.880 6.950 1.040 ;
        RECT  5.950 1.530 6.160 1.690 ;
        RECT  5.340 1.520 5.400 1.760 ;
        RECT  3.600 1.680 3.760 2.040 ;
        RECT  3.480 0.470 3.640 0.790 ;
        RECT  4.600 1.640 5.030 1.800 ;
        RECT  3.930 1.660 4.190 1.800 ;
        RECT  2.440 0.780 2.600 1.950 ;
        RECT  2.060 1.620 2.160 1.780 ;
        RECT  1.080 1.640 1.820 1.800 ;
        RECT  0.060 1.640 0.650 1.800 ;
    END
END SDFXD2

MACRO SDFXD4
    CLASS CORE ;
    FOREIGN SDFXD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.270 3.110 1.795 ;
        RECT  3.110 1.270 3.150 1.510 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.380 3.930 1.540 ;
        RECT  3.930 1.005 4.070 1.540 ;
        END
    END SE
    PIN SA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END SA
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.150 1.650 11.470 2.030 ;
        RECT  11.150 0.490 11.470 0.870 ;
        RECT  11.470 0.490 11.890 2.030 ;
        RECT  11.890 1.650 12.060 2.030 ;
        RECT  11.890 0.490 12.060 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.750 1.600 10.190 1.760 ;
        RECT  9.750 0.760 10.190 0.920 ;
        RECT  10.190 0.760 10.610 1.760 ;
        RECT  10.610 1.600 10.700 1.760 ;
        RECT  10.610 0.760 10.700 0.920 ;
        END
    END Q
    PIN DB
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.110 1.370 1.330 ;
        RECT  1.370 1.005 1.510 1.515 ;
        END
    END DB
    PIN DA
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.970 1.050 1.050 1.270 ;
        RECT  1.050 1.005 1.190 1.515 ;
        END
    END DA
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 4.710 1.515 ;
        RECT  4.710 1.050 4.900 1.270 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.340 ;
        RECT  0.670 -0.300 2.800 0.300 ;
        RECT  2.800 -0.300 3.020 0.760 ;
        RECT  3.020 -0.300 6.540 0.300 ;
        RECT  6.540 -0.300 6.760 0.760 ;
        RECT  6.760 -0.300 12.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.800 2.820 ;
        RECT  2.800 1.920 3.020 2.820 ;
        RECT  3.020 2.220 6.520 2.820 ;
        RECT  6.520 2.030 6.740 2.820 ;
        RECT  6.740 2.220 12.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.630 0.750 1.750 1.050 ;
        RECT  0.810 0.750 1.630 0.870 ;
        RECT  0.650 0.470 0.810 1.800 ;
        RECT  0.060 0.470 0.650 0.630 ;
        RECT  1.990 1.190 2.040 1.350 ;
        RECT  1.940 0.470 1.990 1.350 ;
        RECT  1.870 0.470 1.940 1.800 ;
        RECT  1.070 0.470 1.870 0.630 ;
        RECT  1.820 1.190 1.870 1.800 ;
        RECT  2.280 0.470 2.560 0.630 ;
        RECT  2.160 0.470 2.280 1.780 ;
        RECT  2.110 0.470 2.160 0.690 ;
        RECT  3.460 0.910 3.620 1.560 ;
        RECT  2.600 0.910 3.460 1.070 ;
        RECT  4.190 0.710 4.310 1.800 ;
        RECT  3.830 0.710 4.190 0.870 ;
        RECT  5.150 1.050 5.280 1.270 ;
        RECT  5.030 0.710 5.150 1.800 ;
        RECT  4.500 0.710 5.030 0.870 ;
        RECT  5.520 0.420 5.760 0.590 ;
        RECT  3.640 0.470 5.520 0.590 ;
        RECT  5.580 1.920 5.820 2.080 ;
        RECT  3.760 1.920 5.580 2.040 ;
        RECT  5.520 1.120 6.040 1.280 ;
        RECT  5.400 0.710 5.520 1.760 ;
        RECT  5.300 0.710 5.400 0.930 ;
        RECT  6.830 1.170 6.880 1.410 ;
        RECT  6.710 1.170 6.830 1.690 ;
        RECT  6.280 1.570 6.710 1.690 ;
        RECT  6.160 0.610 6.280 1.690 ;
        RECT  5.890 0.610 6.160 0.770 ;
        RECT  7.000 0.530 7.120 1.930 ;
        RECT  6.950 0.530 7.000 1.040 ;
        RECT  6.950 1.690 7.000 1.930 ;
        RECT  8.960 1.050 9.120 1.480 ;
        RECT  7.490 1.360 8.960 1.480 ;
        RECT  9.505 1.080 9.880 1.240 ;
        RECT  9.385 0.810 9.505 1.810 ;
        RECT  9.300 0.810 9.385 0.930 ;
        RECT  9.060 1.650 9.385 1.810 ;
        RECT  9.080 0.710 9.300 0.930 ;
        RECT  8.660 0.810 9.080 0.930 ;
        RECT  8.540 0.810 8.660 1.240 ;
        RECT  10.980 1.080 11.255 1.240 ;
        RECT  10.860 0.470 10.980 2.050 ;
        RECT  8.610 0.470 10.860 0.590 ;
        RECT  8.580 1.930 10.860 2.050 ;
        RECT  7.870 0.470 8.610 0.630 ;
        RECT  8.360 1.630 8.580 2.050 ;
        RECT  7.660 1.720 8.360 1.880 ;
        RECT  7.710 0.470 7.870 0.805 ;
        RECT  8.420 1.080 8.540 1.240 ;
        RECT  7.330 0.545 7.490 1.930 ;
        RECT  6.410 0.880 6.950 1.040 ;
        RECT  5.950 1.530 6.160 1.690 ;
        RECT  5.340 1.520 5.400 1.760 ;
        RECT  3.600 1.680 3.760 2.040 ;
        RECT  3.480 0.470 3.640 0.790 ;
        RECT  4.600 1.640 5.030 1.800 ;
        RECT  3.930 1.660 4.190 1.800 ;
        RECT  2.440 0.780 2.600 1.950 ;
        RECT  2.060 1.620 2.160 1.780 ;
        RECT  1.080 1.640 1.820 1.800 ;
        RECT  0.060 1.640 0.650 1.800 ;
        LAYER M1 ;
        RECT  11.150 0.490 11.255 0.870 ;
        RECT  9.750 1.600 9.975 1.760 ;
        RECT  9.750 0.760 9.975 0.920 ;
        RECT  11.150 1.650 11.255 2.030 ;
    END
END SDFXD4

MACRO SEDF4CQD1
    CLASS CORE ;
    FOREIGN SEDF4CQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.160 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.070 1.610 11.290 1.770 ;
        RECT  11.070 0.750 11.290 0.910 ;
        RECT  11.290 0.750 11.430 1.770 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.790 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 9.050 0.300 ;
        RECT  9.050 -0.300 9.210 0.770 ;
        RECT  9.210 -0.300 11.470 0.300 ;
        RECT  11.470 -0.300 11.690 0.350 ;
        RECT  11.690 -0.300 12.160 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.820 2.820 ;
        RECT  5.820 2.180 6.040 2.820 ;
        RECT  6.040 2.220 8.950 2.820 ;
        RECT  8.950 2.050 9.170 2.820 ;
        RECT  9.170 2.220 10.430 2.820 ;
        RECT  10.430 2.170 10.650 2.820 ;
        RECT  10.650 2.220 11.470 2.820 ;
        RECT  11.470 2.170 11.690 2.820 ;
        RECT  11.690 2.220 12.160 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.910 0.950 3.030 2.050 ;
        RECT  3.030 0.950 3.170 1.090 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  4.630 1.930 8.700 2.050 ;
        RECT  8.700 1.810 8.820 2.050 ;
        RECT  8.820 1.810 9.395 1.930 ;
        RECT  9.395 1.810 9.515 2.050 ;
        RECT  9.515 1.930 11.900 2.050 ;
        RECT  11.900 0.680 12.060 2.050 ;
        RECT  10.270 0.800 10.830 0.960 ;
        RECT  10.740 0.420 10.830 0.590 ;
        RECT  10.830 0.420 10.950 1.800 ;
        RECT  10.950 0.420 10.980 0.590 ;
        RECT  10.980 0.470 11.580 0.590 ;
        RECT  11.580 0.470 11.740 1.300 ;
        RECT  10.020 0.420 10.140 1.270 ;
        RECT  9.710 1.670 10.400 1.810 ;
        RECT  10.140 1.140 10.400 1.270 ;
        RECT  10.400 1.140 10.520 1.810 ;
        RECT  10.520 1.140 10.710 1.360 ;
        RECT  9.850 1.390 10.160 1.550 ;
        RECT  8.980 1.440 9.460 1.600 ;
        RECT  9.430 0.530 9.460 0.770 ;
        RECT  9.460 0.530 9.580 1.600 ;
        RECT  8.350 0.670 8.450 0.830 ;
        RECT  8.450 0.670 8.570 1.600 ;
        RECT  8.570 0.670 8.590 1.010 ;
        RECT  8.590 0.890 9.170 1.010 ;
        RECT  9.170 0.890 9.330 1.280 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.260 1.690 7.950 1.810 ;
        RECT  7.950 1.380 8.020 1.810 ;
        RECT  5.510 0.470 8.020 0.590 ;
        RECT  8.020 0.470 8.110 1.810 ;
        RECT  8.110 0.470 8.180 1.500 ;
        RECT  7.545 0.720 7.665 1.570 ;
        RECT  7.665 0.720 7.705 1.220 ;
        RECT  7.705 1.060 7.900 1.220 ;
        RECT  6.630 0.750 6.760 0.910 ;
        RECT  6.760 0.750 6.880 1.570 ;
        RECT  6.880 1.080 7.425 1.240 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.270 ;
        RECT  6.510 1.050 6.640 1.270 ;
        RECT  5.560 0.740 5.940 0.880 ;
        RECT  5.940 0.740 6.060 1.570 ;
        RECT  6.060 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.240 1.600 ;
        RECT  1.240 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  10.710 1.640 10.830 1.800 ;
        RECT  9.760 0.420 10.020 0.560 ;
        RECT  9.700 0.790 9.850 1.550 ;
        RECT  8.820 1.140 8.980 1.600 ;
        RECT  8.330 1.380 8.450 1.600 ;
        RECT  7.330 1.410 7.545 1.570 ;
        RECT  6.600 1.410 6.760 1.570 ;
        RECT  6.190 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.940 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  2.670 1.620 2.910 1.780 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDF4CQD1

MACRO SEDF4CQD2
    CLASS CORE ;
    FOREIGN SEDF4CQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.370 1.610 11.610 1.770 ;
        RECT  11.390 0.750 11.610 0.910 ;
        RECT  11.610 0.750 11.750 1.770 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.790 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 9.050 0.300 ;
        RECT  9.050 -0.300 9.210 0.770 ;
        RECT  9.210 -0.300 11.810 0.300 ;
        RECT  11.810 -0.300 12.030 0.340 ;
        RECT  12.030 -0.300 12.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.820 2.820 ;
        RECT  5.820 2.180 6.040 2.820 ;
        RECT  6.040 2.220 8.950 2.820 ;
        RECT  8.950 2.050 9.170 2.820 ;
        RECT  9.170 2.220 10.430 2.820 ;
        RECT  10.430 2.190 10.650 2.820 ;
        RECT  10.650 2.220 10.970 2.820 ;
        RECT  10.970 2.180 11.190 2.820 ;
        RECT  11.190 2.220 11.790 2.820 ;
        RECT  11.790 2.170 12.010 2.820 ;
        RECT  12.010 2.220 12.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  4.630 1.930 8.700 2.050 ;
        RECT  8.700 1.810 8.820 2.050 ;
        RECT  8.820 1.810 9.395 1.930 ;
        RECT  9.395 1.810 9.515 2.050 ;
        RECT  9.515 1.930 12.220 2.050 ;
        RECT  12.220 0.680 12.380 2.050 ;
        RECT  10.270 0.800 10.830 0.960 ;
        RECT  10.740 0.420 10.830 0.590 ;
        RECT  10.830 0.420 10.950 1.800 ;
        RECT  10.950 0.420 10.980 0.590 ;
        RECT  10.980 0.470 11.940 0.590 ;
        RECT  11.940 0.470 12.100 1.300 ;
        RECT  10.020 0.420 10.140 1.270 ;
        RECT  9.710 1.670 10.400 1.810 ;
        RECT  10.140 1.140 10.400 1.270 ;
        RECT  10.400 1.140 10.520 1.810 ;
        RECT  10.520 1.140 10.710 1.360 ;
        RECT  9.850 1.390 10.160 1.550 ;
        RECT  8.980 1.440 9.460 1.600 ;
        RECT  9.430 0.530 9.460 0.770 ;
        RECT  9.460 0.530 9.580 1.600 ;
        RECT  8.350 0.670 8.450 0.830 ;
        RECT  8.450 0.670 8.570 1.600 ;
        RECT  8.570 0.670 8.590 1.010 ;
        RECT  8.590 0.890 9.170 1.010 ;
        RECT  9.170 0.890 9.330 1.280 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.260 1.690 7.950 1.810 ;
        RECT  7.950 1.380 8.020 1.810 ;
        RECT  5.510 0.470 8.020 0.590 ;
        RECT  8.020 0.470 8.110 1.810 ;
        RECT  8.110 0.470 8.180 1.500 ;
        RECT  7.545 0.720 7.665 1.570 ;
        RECT  7.665 0.720 7.705 1.220 ;
        RECT  7.705 1.060 7.900 1.220 ;
        RECT  6.630 0.750 6.760 0.910 ;
        RECT  6.760 0.750 6.880 1.570 ;
        RECT  6.880 1.080 7.425 1.240 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.270 ;
        RECT  6.510 1.050 6.640 1.270 ;
        RECT  5.560 0.740 5.940 0.880 ;
        RECT  5.940 0.740 6.060 1.570 ;
        RECT  6.060 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.240 1.600 ;
        RECT  1.240 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.030 0.950 3.170 1.090 ;
        RECT  2.910 0.950 3.030 2.050 ;
        RECT  10.710 1.640 10.830 1.800 ;
        RECT  9.760 0.420 10.020 0.560 ;
        RECT  9.700 0.790 9.850 1.550 ;
        RECT  8.820 1.140 8.980 1.600 ;
        RECT  8.330 1.380 8.450 1.600 ;
        RECT  7.330 1.410 7.545 1.570 ;
        RECT  6.600 1.410 6.760 1.570 ;
        RECT  6.190 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.940 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  2.670 1.620 2.910 1.780 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDF4CQD2

MACRO SEDF4CQD4
    CLASS CORE ;
    FOREIGN SEDF4CQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.630 1.610 12.750 1.770 ;
        RECT  12.670 0.750 12.750 0.910 ;
        RECT  12.750 0.750 13.170 1.770 ;
        RECT  13.170 1.610 13.580 1.770 ;
        RECT  13.170 0.750 13.620 0.910 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.790 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 9.050 0.300 ;
        RECT  9.050 -0.300 9.210 0.770 ;
        RECT  9.210 -0.300 9.840 0.300 ;
        RECT  9.840 -0.300 10.060 0.485 ;
        RECT  10.060 -0.300 13.780 0.300 ;
        RECT  13.780 -0.300 14.000 0.340 ;
        RECT  14.000 -0.300 14.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.820 2.820 ;
        RECT  5.820 2.180 6.040 2.820 ;
        RECT  6.040 2.220 8.950 2.820 ;
        RECT  8.950 2.050 9.170 2.820 ;
        RECT  9.170 2.220 9.750 2.820 ;
        RECT  9.750 2.050 9.970 2.820 ;
        RECT  9.970 2.220 11.650 2.820 ;
        RECT  11.650 2.180 11.870 2.820 ;
        RECT  11.870 2.220 12.250 2.820 ;
        RECT  12.250 2.180 12.470 2.820 ;
        RECT  12.470 2.220 13.740 2.820 ;
        RECT  13.740 2.180 13.960 2.820 ;
        RECT  13.960 2.220 14.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.740 1.140 11.930 1.360 ;
        RECT  11.080 1.400 11.380 1.550 ;
        RECT  8.980 1.440 9.460 1.600 ;
        RECT  9.430 0.530 9.460 0.770 ;
        RECT  9.460 0.530 9.580 1.600 ;
        RECT  9.580 1.065 10.570 1.185 ;
        RECT  10.570 0.740 10.690 1.550 ;
        RECT  10.690 1.410 10.810 1.550 ;
        RECT  10.690 0.740 10.820 0.900 ;
        RECT  8.350 0.670 8.450 0.830 ;
        RECT  8.450 0.670 8.570 1.600 ;
        RECT  8.570 0.670 8.590 1.010 ;
        RECT  8.590 0.890 9.170 1.010 ;
        RECT  9.170 0.890 9.330 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.260 1.690 7.950 1.810 ;
        RECT  7.950 1.380 8.020 1.810 ;
        RECT  5.510 0.470 8.020 0.590 ;
        RECT  8.020 0.470 8.110 1.810 ;
        RECT  8.110 0.470 8.180 1.500 ;
        RECT  7.545 0.720 7.665 1.570 ;
        RECT  7.665 0.720 7.705 1.220 ;
        RECT  7.705 1.060 7.900 1.220 ;
        RECT  6.630 0.750 6.760 0.910 ;
        RECT  6.760 0.750 6.880 1.570 ;
        RECT  6.880 1.080 7.425 1.240 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.270 ;
        RECT  6.510 1.050 6.640 1.270 ;
        RECT  5.560 0.740 5.940 0.880 ;
        RECT  5.940 0.740 6.060 1.570 ;
        RECT  6.060 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.240 1.600 ;
        RECT  1.240 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  11.620 1.140 11.740 1.810 ;
        RECT  11.360 1.140 11.620 1.270 ;
        RECT  10.450 1.670 11.620 1.810 ;
        RECT  11.240 0.470 11.360 1.270 ;
        RECT  10.420 0.470 11.240 0.610 ;
        RECT  10.330 1.465 10.450 1.810 ;
        RECT  10.180 0.470 10.420 0.630 ;
        RECT  13.880 0.470 14.020 1.300 ;
        RECT  12.200 0.470 13.880 0.590 ;
        RECT  12.170 0.420 12.200 0.590 ;
        RECT  12.050 0.420 12.170 1.800 ;
        RECT  11.960 0.420 12.050 0.590 ;
        RECT  11.490 0.800 12.050 0.960 ;
        RECT  14.140 0.680 14.300 2.050 ;
        RECT  10.210 1.930 14.140 2.050 ;
        RECT  10.090 1.810 10.210 2.050 ;
        RECT  8.820 1.810 10.090 1.930 ;
        RECT  8.700 1.810 8.820 2.050 ;
        RECT  4.630 1.930 8.700 2.050 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.030 0.950 3.170 1.090 ;
        RECT  2.910 0.950 3.030 2.050 ;
        RECT  11.930 1.640 12.050 1.800 ;
        RECT  10.170 1.465 10.330 1.625 ;
        RECT  10.940 0.810 11.080 1.550 ;
        RECT  8.820 1.140 8.980 1.600 ;
        RECT  8.330 1.380 8.450 1.600 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  7.330 1.410 7.545 1.570 ;
        RECT  6.600 1.410 6.760 1.570 ;
        RECT  6.190 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.940 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  2.670 1.620 2.910 1.780 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
        LAYER M1 ;
        RECT  13.385 0.750 13.620 0.910 ;
        RECT  13.385 1.610 13.580 1.770 ;
    END
END SEDF4CQD4

MACRO SEDFCND1
    CLASS CORE ;
    FOREIGN SEDFCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.230 1.940 11.260 2.100 ;
        RECT  11.260 1.390 11.290 2.100 ;
        RECT  11.260 0.420 11.290 0.920 ;
        RECT  11.290 0.420 11.420 2.100 ;
        RECT  11.420 0.800 11.430 1.515 ;
        RECT  11.420 1.940 11.450 2.100 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.445 1.600 10.650 1.760 ;
        RECT  10.515 0.710 10.650 0.930 ;
        RECT  10.650 0.710 10.655 1.760 ;
        RECT  10.655 0.810 10.790 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.970 1.140 10.010 1.360 ;
        RECT  10.010 1.140 10.150 1.795 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 11.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 4.540 2.820 ;
        RECT  4.540 2.180 4.760 2.820 ;
        RECT  4.760 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 10.050 2.820 ;
        RECT  10.050 2.180 10.270 2.820 ;
        RECT  10.270 2.220 11.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.920 1.410 9.050 1.570 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.270 1.930 10.990 2.050 ;
        RECT  9.850 0.470 10.990 0.590 ;
        RECT  10.990 0.470 11.110 2.050 ;
        RECT  11.110 1.050 11.170 1.270 ;
        RECT  9.180 0.900 9.300 1.270 ;
        RECT  9.620 1.670 9.730 1.810 ;
        RECT  9.300 0.900 9.730 1.020 ;
        RECT  9.730 0.900 9.850 1.810 ;
        RECT  9.850 1.670 9.860 1.810 ;
        RECT  9.850 0.900 10.040 1.020 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  10.260 0.900 10.270 1.020 ;
        RECT  10.270 0.900 10.390 1.270 ;
        RECT  10.390 1.050 10.530 1.270 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.620 1.690 9.180 1.810 ;
        RECT  9.180 1.420 9.300 1.810 ;
        RECT  9.300 1.420 9.470 1.540 ;
        RECT  9.470 1.140 9.610 1.540 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.860 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.020 2.150 1.180 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.110 9.180 1.270 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
    END
END SEDFCND1

MACRO SEDFCND2
    CLASS CORE ;
    FOREIGN SEDFCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.790 1.940 11.820 2.100 ;
        RECT  11.820 1.390 11.980 2.100 ;
        RECT  11.820 0.420 11.980 0.920 ;
        RECT  11.980 1.940 12.010 2.100 ;
        RECT  11.980 1.390 12.250 1.515 ;
        RECT  11.980 0.800 12.250 0.920 ;
        RECT  12.250 0.800 12.390 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.150 1.570 11.290 1.810 ;
        RECT  11.150 0.710 11.290 0.950 ;
        RECT  11.290 0.830 11.430 1.690 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.330 1.285 10.545 1.515 ;
        RECT  10.545 1.105 10.710 1.515 ;
        RECT  10.710 1.285 10.790 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 10.690 0.300 ;
        RECT  10.690 -0.300 10.910 0.340 ;
        RECT  10.910 -0.300 12.480 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 4.540 2.820 ;
        RECT  4.540 2.180 4.760 2.820 ;
        RECT  4.760 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 12.480 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  11.550 0.470 11.670 2.050 ;
        RECT  11.670 1.080 11.900 1.240 ;
        RECT  9.640 0.900 9.760 1.570 ;
        RECT  9.760 1.430 9.860 1.570 ;
        RECT  9.760 0.900 10.040 1.020 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  10.325 1.635 10.910 1.795 ;
        RECT  10.260 0.710 10.910 0.830 ;
        RECT  10.910 0.710 11.030 1.795 ;
        RECT  11.030 1.050 11.050 1.270 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.620 1.690 9.980 1.810 ;
        RECT  9.980 1.140 10.140 1.810 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.860 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.020 2.150 1.180 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  9.850 0.470 11.550 0.590 ;
        RECT  8.270 1.930 11.550 2.050 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  8.920 1.410 9.070 1.570 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.110 9.640 1.270 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
    END
END SEDFCND2

MACRO SEDFCND4
    CLASS CORE ;
    FOREIGN SEDFCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  13.070 1.650 13.390 2.030 ;
        RECT  13.070 0.490 13.390 0.870 ;
        RECT  13.390 0.490 13.810 2.030 ;
        RECT  13.810 1.650 13.980 2.030 ;
        RECT  13.810 0.490 13.980 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.670 1.600 11.790 1.760 ;
        RECT  11.670 0.760 11.790 0.920 ;
        RECT  11.790 0.760 12.210 1.760 ;
        RECT  12.210 1.600 12.620 1.760 ;
        RECT  12.210 0.760 12.620 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.545 1.125 10.650 1.360 ;
        RECT  10.650 1.005 10.790 1.515 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 14.400 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 14.400 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.830 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.080 2.150 1.240 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  10.035 1.140 10.195 1.810 ;
        RECT  8.620 1.690 10.035 1.810 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  11.260 0.710 11.420 1.800 ;
        RECT  10.260 0.710 11.260 0.830 ;
        RECT  10.320 1.640 11.260 1.800 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  9.760 0.900 10.040 1.020 ;
        RECT  9.760 1.430 9.880 1.570 ;
        RECT  9.640 0.900 9.760 1.570 ;
        RECT  12.900 1.080 13.175 1.240 ;
        RECT  12.780 0.470 12.900 2.050 ;
        RECT  9.850 0.470 12.780 0.590 ;
        RECT  8.270 1.930 12.780 2.050 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  8.920 1.410 9.070 1.570 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.030 9.640 1.190 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
        LAYER M1 ;
        RECT  13.070 1.650 13.175 2.030 ;
        RECT  13.070 0.490 13.175 0.870 ;
        RECT  12.425 1.600 12.620 1.760 ;
        RECT  12.425 0.760 12.620 0.920 ;
    END
END SEDFCND4

MACRO SEDFCNQD1
    CLASS CORE ;
    FOREIGN SEDFCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.445 1.600 10.650 1.760 ;
        RECT  10.515 0.710 10.650 0.930 ;
        RECT  10.650 0.710 10.655 1.760 ;
        RECT  10.655 0.810 10.790 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.970 1.140 10.010 1.360 ;
        RECT  10.010 1.140 10.150 1.795 ;
        END
    END CDN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 4.540 2.820 ;
        RECT  4.540 2.180 4.760 2.820 ;
        RECT  4.760 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 10.050 2.820 ;
        RECT  10.050 2.180 10.270 2.820 ;
        RECT  10.270 2.220 10.860 2.820 ;
        RECT  10.860 2.180 11.080 2.820 ;
        RECT  11.080 2.220 11.200 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 10.860 0.300 ;
        RECT  10.860 -0.300 11.080 0.340 ;
        RECT  11.080 -0.300 11.200 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  9.180 0.900 9.300 1.270 ;
        RECT  9.620 1.670 9.730 1.810 ;
        RECT  9.300 0.900 9.730 1.020 ;
        RECT  9.730 0.900 9.850 1.810 ;
        RECT  9.850 1.670 9.860 1.810 ;
        RECT  9.850 0.900 10.040 1.020 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  10.260 0.900 10.270 1.020 ;
        RECT  10.270 0.900 10.390 1.270 ;
        RECT  10.390 1.050 10.530 1.270 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.620 1.690 9.180 1.810 ;
        RECT  9.180 1.420 9.300 1.810 ;
        RECT  9.300 1.420 9.470 1.540 ;
        RECT  9.470 1.140 9.610 1.540 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.860 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.020 2.150 1.180 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  10.990 0.470 11.110 2.050 ;
        RECT  9.850 0.470 10.990 0.590 ;
        RECT  8.270 1.930 10.990 2.050 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  8.920 1.410 9.050 1.570 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.110 9.180 1.270 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
    END
END SEDFCNQD1

MACRO SEDFCNQD2
    CLASS CORE ;
    FOREIGN SEDFCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.150 1.570 11.290 1.810 ;
        RECT  11.150 0.710 11.290 0.950 ;
        RECT  11.290 0.830 11.430 1.690 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.330 1.285 10.545 1.515 ;
        RECT  10.545 1.105 10.710 1.515 ;
        RECT  10.710 1.285 10.790 1.515 ;
        END
    END CDN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 4.540 2.820 ;
        RECT  4.540 2.180 4.760 2.820 ;
        RECT  4.760 2.220 5.080 2.820 ;
        RECT  5.080 2.180 5.300 2.820 ;
        RECT  5.300 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 11.500 2.820 ;
        RECT  11.500 2.180 11.720 2.820 ;
        RECT  11.720 2.220 11.840 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 4.450 0.300 ;
        RECT  4.450 -0.300 4.670 0.340 ;
        RECT  4.670 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 10.690 0.300 ;
        RECT  10.690 -0.300 10.910 0.340 ;
        RECT  10.910 -0.300 11.500 0.300 ;
        RECT  11.500 -0.300 11.720 0.340 ;
        RECT  11.720 -0.300 11.840 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  9.640 0.900 9.760 1.570 ;
        RECT  9.760 1.430 9.860 1.570 ;
        RECT  9.760 0.900 10.040 1.020 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  10.325 1.635 10.910 1.795 ;
        RECT  10.260 0.710 10.910 0.830 ;
        RECT  10.910 0.710 11.030 1.795 ;
        RECT  11.030 1.050 11.050 1.270 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.620 1.690 9.980 1.810 ;
        RECT  9.980 1.140 10.140 1.810 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.830 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.020 2.150 1.180 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  11.550 0.470 11.670 2.050 ;
        RECT  9.850 0.470 11.550 0.590 ;
        RECT  8.270 1.930 11.550 2.050 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  8.920 1.410 9.070 1.570 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.110 9.640 1.270 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
    END
END SEDFCNQD2

MACRO SEDFCNQD4
    CLASS CORE ;
    FOREIGN SEDFCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.480 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.285 3.430 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.070 1.515 ;
        RECT  4.070 1.060 4.190 1.230 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.150 1.600 11.470 1.760 ;
        RECT  11.150 0.760 11.470 0.920 ;
        RECT  11.470 0.760 11.890 1.760 ;
        RECT  11.890 1.600 12.080 1.760 ;
        RECT  11.890 0.760 12.080 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.235 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.730 0.725 1.190 0.955 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.005 5.030 1.235 ;
        END
    END CP
    PIN CDN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  10.545 1.125 10.650 1.360 ;
        RECT  10.650 1.005 10.790 1.515 ;
        END
    END CDN
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.440 2.820 ;
        RECT  0.440 1.690 0.660 2.820 ;
        RECT  0.660 2.220 1.700 2.820 ;
        RECT  1.700 1.690 1.920 2.820 ;
        RECT  1.920 2.220 3.070 2.820 ;
        RECT  3.070 1.880 3.290 2.820 ;
        RECT  3.290 2.220 6.970 2.820 ;
        RECT  6.970 2.060 7.190 2.820 ;
        RECT  7.190 2.220 7.640 2.820 ;
        RECT  7.640 2.060 7.860 2.820 ;
        RECT  7.860 2.220 9.245 2.820 ;
        RECT  9.245 2.180 9.465 2.820 ;
        RECT  9.465 2.220 10.750 2.820 ;
        RECT  10.750 2.180 10.970 2.820 ;
        RECT  10.970 2.220 12.480 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.340 ;
        RECT  1.950 -0.300 2.890 0.300 ;
        RECT  2.890 -0.300 3.110 0.920 ;
        RECT  3.110 -0.300 4.440 0.300 ;
        RECT  4.440 -0.300 4.660 0.340 ;
        RECT  4.660 -0.300 7.140 0.300 ;
        RECT  7.140 -0.300 7.360 0.490 ;
        RECT  7.360 -0.300 9.390 0.300 ;
        RECT  9.390 -0.300 9.610 0.480 ;
        RECT  9.610 -0.300 10.750 0.300 ;
        RECT  10.750 -0.300 10.970 0.340 ;
        RECT  10.970 -0.300 12.480 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  10.320 1.640 10.910 1.800 ;
        RECT  10.260 0.710 10.910 0.830 ;
        RECT  10.910 0.710 11.030 1.800 ;
        RECT  8.270 1.140 8.460 1.260 ;
        RECT  8.460 1.140 8.620 1.810 ;
        RECT  8.620 1.690 10.035 1.810 ;
        RECT  10.035 1.140 10.195 1.810 ;
        RECT  6.960 1.320 7.720 1.440 ;
        RECT  7.720 0.710 7.880 1.645 ;
        RECT  7.880 1.485 8.290 1.645 ;
        RECT  6.590 0.730 7.480 0.850 ;
        RECT  7.480 0.470 7.600 0.850 ;
        RECT  7.600 0.470 7.960 0.590 ;
        RECT  7.960 0.430 8.180 0.590 ;
        RECT  6.250 0.420 6.310 1.610 ;
        RECT  6.310 1.040 6.410 1.610 ;
        RECT  6.410 1.040 7.380 1.160 ;
        RECT  7.380 1.040 7.600 1.200 ;
        RECT  6.540 1.560 7.460 1.700 ;
        RECT  3.940 1.690 6.070 1.810 ;
        RECT  3.810 0.470 5.740 0.590 ;
        RECT  5.740 0.430 5.980 0.590 ;
        RECT  5.390 0.710 5.660 0.830 ;
        RECT  5.660 0.710 5.820 1.570 ;
        RECT  4.680 0.710 5.150 0.830 ;
        RECT  5.150 0.710 5.270 1.570 ;
        RECT  5.270 0.985 5.490 1.145 ;
        RECT  4.030 0.710 4.330 0.830 ;
        RECT  4.330 0.710 4.450 1.570 ;
        RECT  2.700 1.040 3.600 1.160 ;
        RECT  3.600 1.040 3.760 1.325 ;
        RECT  2.110 0.470 2.270 0.630 ;
        RECT  2.270 0.470 2.390 1.590 ;
        RECT  2.390 0.470 2.620 0.610 ;
        RECT  1.050 0.440 1.290 0.600 ;
        RECT  1.260 1.450 1.540 1.570 ;
        RECT  1.290 0.480 1.540 0.600 ;
        RECT  1.540 0.480 1.660 1.570 ;
        RECT  1.660 1.080 2.150 1.240 ;
        RECT  0.060 0.430 0.280 0.590 ;
        RECT  0.250 1.430 0.410 1.550 ;
        RECT  0.280 0.470 0.410 0.590 ;
        RECT  0.410 0.470 0.530 1.550 ;
        RECT  0.530 1.100 1.420 1.260 ;
        RECT  10.040 0.710 10.260 1.020 ;
        RECT  9.760 0.900 10.040 1.020 ;
        RECT  9.760 1.430 9.880 1.570 ;
        RECT  9.640 0.900 9.760 1.570 ;
        RECT  12.240 0.470 12.360 2.050 ;
        RECT  9.850 0.470 12.240 0.590 ;
        RECT  8.270 1.930 12.240 2.050 ;
        RECT  9.730 0.470 9.850 0.780 ;
        RECT  8.920 0.640 9.730 0.780 ;
        RECT  8.920 1.410 9.070 1.570 ;
        RECT  8.800 0.640 8.920 1.570 ;
        RECT  8.560 0.780 8.800 0.940 ;
        RECT  8.150 1.820 8.270 2.050 ;
        RECT  6.330 1.820 8.150 1.940 ;
        RECT  6.210 1.820 6.330 2.050 ;
        RECT  3.560 1.930 6.210 2.050 ;
        RECT  3.440 1.640 3.560 2.050 ;
        RECT  2.950 1.640 3.440 1.760 ;
        RECT  2.830 1.640 2.950 2.050 ;
        RECT  2.610 1.930 2.830 2.050 ;
        RECT  9.060 1.030 9.640 1.190 ;
        RECT  2.390 1.930 2.610 2.100 ;
        RECT  8.110 0.720 8.270 1.260 ;
        RECT  6.720 1.280 6.960 1.440 ;
        RECT  6.430 0.420 6.590 0.850 ;
        RECT  6.150 0.420 6.250 1.160 ;
        RECT  3.700 1.650 3.940 1.810 ;
        RECT  3.590 0.470 3.810 0.730 ;
        RECT  5.460 1.410 5.660 1.570 ;
        RECT  4.770 1.410 5.150 1.570 ;
        RECT  4.190 1.350 4.330 1.570 ;
        RECT  2.540 0.730 2.700 1.810 ;
        RECT  2.110 1.470 2.270 1.950 ;
        RECT  1.100 1.450 1.260 1.900 ;
        RECT  0.090 1.430 0.250 1.900 ;
        LAYER M1 ;
        RECT  11.150 1.600 11.255 1.760 ;
        RECT  11.150 0.760 11.255 0.920 ;
    END
END SEDFCNQD4

MACRO SEDFD1
    CLASS CORE ;
    FOREIGN SEDFD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.190 1.940 11.220 2.100 ;
        RECT  11.220 1.390 11.290 2.100 ;
        RECT  11.220 0.420 11.290 0.920 ;
        RECT  11.290 0.420 11.390 2.100 ;
        RECT  11.390 1.940 11.410 2.100 ;
        RECT  11.390 0.800 11.430 1.515 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.660 1.580 9.690 1.800 ;
        RECT  9.660 0.720 9.690 0.940 ;
        RECT  9.690 0.720 9.830 1.800 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.350 ;
        RECT  6.110 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 10.030 0.300 ;
        RECT  10.030 -0.300 10.250 0.340 ;
        RECT  10.250 -0.300 10.790 0.300 ;
        RECT  10.790 -0.300 11.010 0.340 ;
        RECT  11.010 -0.300 11.520 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.730 2.820 ;
        RECT  5.730 2.170 5.950 2.820 ;
        RECT  5.950 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 8.990 2.820 ;
        RECT  8.990 2.170 9.210 2.820 ;
        RECT  9.210 2.220 10.030 2.820 ;
        RECT  10.030 2.180 10.250 2.820 ;
        RECT  10.250 2.220 10.790 2.820 ;
        RECT  10.790 2.180 11.010 2.820 ;
        RECT  11.010 2.220 11.520 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  7.380 1.810 7.955 1.930 ;
        RECT  7.955 1.810 8.075 2.050 ;
        RECT  8.075 1.930 10.530 2.050 ;
        RECT  10.410 1.520 10.530 1.680 ;
        RECT  10.410 0.730 10.530 0.890 ;
        RECT  10.530 0.730 10.650 2.050 ;
        RECT  8.830 0.800 9.390 0.960 ;
        RECT  9.300 0.420 9.390 0.590 ;
        RECT  9.390 0.420 9.510 1.800 ;
        RECT  9.510 0.420 9.540 0.590 ;
        RECT  9.540 0.470 10.150 0.590 ;
        RECT  10.150 0.470 10.270 1.280 ;
        RECT  10.270 1.060 10.410 1.280 ;
        RECT  8.580 0.420 8.700 1.270 ;
        RECT  8.270 1.670 8.960 1.810 ;
        RECT  8.700 1.140 8.960 1.270 ;
        RECT  8.960 1.140 9.080 1.810 ;
        RECT  9.080 1.140 9.270 1.360 ;
        RECT  8.410 1.390 8.720 1.550 ;
        RECT  7.540 1.440 8.020 1.600 ;
        RECT  7.990 0.530 8.020 0.770 ;
        RECT  8.020 0.530 8.140 1.600 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.560 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  9.270 1.640 9.390 1.800 ;
        RECT  8.320 0.420 8.580 0.560 ;
        RECT  8.260 0.790 8.410 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDFD1

MACRO SEDFD2
    CLASS CORE ;
    FOREIGN SEDFD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.840 1.610 10.970 1.770 ;
        RECT  10.840 0.750 10.970 0.910 ;
        RECT  10.970 0.750 11.110 1.770 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.010 0.750 10.150 1.770 ;
        RECT  10.150 1.610 10.320 1.770 ;
        RECT  10.150 0.750 10.320 0.910 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.350 ;
        RECT  6.110 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 9.680 0.300 ;
        RECT  9.680 -0.300 9.900 0.340 ;
        RECT  9.900 -0.300 10.470 0.300 ;
        RECT  10.470 -0.300 10.690 0.340 ;
        RECT  10.690 -0.300 11.260 0.300 ;
        RECT  11.260 -0.300 11.480 0.340 ;
        RECT  11.480 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.730 2.820 ;
        RECT  5.730 2.170 5.950 2.820 ;
        RECT  5.950 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 8.990 2.820 ;
        RECT  8.990 2.170 9.210 2.820 ;
        RECT  9.210 2.220 9.680 2.820 ;
        RECT  9.680 2.180 9.900 2.820 ;
        RECT  9.900 2.220 10.470 2.820 ;
        RECT  10.470 2.180 10.690 2.820 ;
        RECT  10.690 2.220 11.260 2.820 ;
        RECT  11.260 2.180 11.480 2.820 ;
        RECT  11.480 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  7.380 1.810 7.955 1.930 ;
        RECT  7.955 1.810 8.075 2.050 ;
        RECT  8.075 1.930 11.580 2.050 ;
        RECT  11.580 0.680 11.740 2.050 ;
        RECT  8.830 0.800 9.390 0.960 ;
        RECT  9.300 0.470 9.390 0.630 ;
        RECT  9.390 0.470 9.510 1.800 ;
        RECT  9.510 0.470 11.280 0.630 ;
        RECT  11.280 0.470 11.440 1.300 ;
        RECT  8.580 0.420 8.700 1.270 ;
        RECT  8.270 1.670 8.960 1.810 ;
        RECT  8.700 1.140 8.960 1.270 ;
        RECT  8.960 1.140 9.080 1.810 ;
        RECT  9.080 1.140 9.270 1.360 ;
        RECT  8.410 1.390 8.720 1.550 ;
        RECT  7.540 1.440 8.020 1.600 ;
        RECT  7.990 0.530 8.020 0.770 ;
        RECT  8.020 0.530 8.140 1.600 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.560 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  9.270 1.640 9.390 1.800 ;
        RECT  8.320 0.420 8.580 0.560 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  8.260 0.790 8.410 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDFD2

MACRO SEDFD4
    CLASS CORE ;
    FOREIGN SEDFD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.390 1.520 12.750 1.680 ;
        RECT  12.390 0.750 12.750 0.910 ;
        RECT  12.750 0.750 13.170 1.680 ;
        RECT  13.170 1.520 13.340 1.680 ;
        RECT  13.170 0.750 13.340 0.910 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.010 1.520 11.150 1.680 ;
        RECT  11.010 0.750 11.150 0.910 ;
        RECT  11.150 0.750 11.570 1.680 ;
        RECT  11.570 1.520 11.960 1.680 ;
        RECT  11.570 0.750 11.960 0.910 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 13.500 0.300 ;
        RECT  13.500 -0.300 13.720 0.340 ;
        RECT  13.720 -0.300 14.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 10.050 2.820 ;
        RECT  10.050 2.170 10.270 2.820 ;
        RECT  10.270 2.220 10.630 2.820 ;
        RECT  10.630 2.170 10.850 2.820 ;
        RECT  10.850 2.220 13.500 2.820 ;
        RECT  13.500 2.180 13.720 2.820 ;
        RECT  13.720 2.220 14.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.400 1.930 13.820 2.050 ;
        RECT  13.820 0.680 13.980 2.050 ;
        RECT  9.890 0.800 10.480 0.960 ;
        RECT  10.360 0.420 10.480 0.590 ;
        RECT  10.480 0.420 10.600 1.680 ;
        RECT  10.600 0.470 13.510 0.590 ;
        RECT  13.510 0.470 13.670 1.300 ;
        RECT  8.660 0.720 8.780 1.810 ;
        RECT  8.780 0.720 8.820 1.410 ;
        RECT  9.380 0.420 9.640 0.560 ;
        RECT  9.640 0.420 9.760 1.290 ;
        RECT  8.780 1.670 10.020 1.810 ;
        RECT  9.760 1.170 10.020 1.290 ;
        RECT  10.020 1.170 10.140 1.810 ;
        RECT  10.140 1.170 10.360 1.330 ;
        RECT  9.470 1.410 9.780 1.550 ;
        RECT  7.540 1.440 8.010 1.600 ;
        RECT  8.010 0.470 8.160 1.600 ;
        RECT  8.970 1.400 9.000 1.550 ;
        RECT  8.160 0.470 9.000 0.590 ;
        RECT  9.000 0.470 9.160 1.550 ;
        RECT  9.160 1.400 9.190 1.550 ;
        RECT  9.160 0.470 9.260 0.630 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.550 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  8.280 1.810 8.400 2.050 ;
        RECT  7.380 1.810 8.280 1.930 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  10.330 1.520 10.480 1.680 ;
        RECT  8.620 1.290 8.660 1.810 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  9.320 0.790 9.470 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
        LAYER M1 ;
        RECT  11.785 0.750 11.960 0.910 ;
        RECT  11.785 1.520 11.960 1.680 ;
        RECT  12.390 0.750 12.535 0.910 ;
        RECT  12.390 1.520 12.535 1.680 ;
    END
END SEDFD4

MACRO SEDFKCND1
    CLASS CORE ;
    FOREIGN SEDFKCND1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.940 1.570 10.970 2.070 ;
        RECT  10.940 0.420 10.970 0.920 ;
        RECT  10.970 0.420 11.100 2.070 ;
        RECT  11.100 0.800 11.110 1.690 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.110 1.600 10.330 1.760 ;
        RECT  10.110 0.710 10.330 0.870 ;
        RECT  10.330 0.710 10.470 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.000 0.300 ;
        RECT  5.000 -0.300 5.220 0.340 ;
        RECT  5.220 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 10.510 0.300 ;
        RECT  10.510 -0.300 10.730 0.340 ;
        RECT  10.730 -0.300 11.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 5.230 2.820 ;
        RECT  5.230 2.180 5.450 2.820 ;
        RECT  5.450 2.220 5.830 2.820 ;
        RECT  5.830 2.180 6.050 2.820 ;
        RECT  6.050 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 9.350 2.820 ;
        RECT  9.350 2.180 9.570 2.820 ;
        RECT  9.570 2.220 10.510 2.820 ;
        RECT  10.510 2.180 10.730 2.820 ;
        RECT  10.730 2.220 11.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  10.810 1.050 10.850 1.270 ;
        RECT  9.290 0.710 9.410 1.240 ;
        RECT  9.730 1.600 9.870 1.760 ;
        RECT  9.410 0.710 9.870 0.870 ;
        RECT  9.870 0.710 9.990 1.760 ;
        RECT  9.990 1.050 10.210 1.270 ;
        RECT  8.330 0.460 8.440 1.740 ;
        RECT  8.440 1.360 8.490 1.740 ;
        RECT  8.490 1.360 9.560 1.480 ;
        RECT  9.560 1.030 9.720 1.480 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.330 1.720 ;
        RECT  3.330 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  10.690 0.470 10.810 2.050 ;
        RECT  9.280 0.470 10.690 0.590 ;
        RECT  8.970 1.930 10.690 2.050 ;
        RECT  9.060 0.430 9.280 0.590 ;
        RECT  8.830 0.470 9.060 0.590 ;
        RECT  8.750 1.630 8.970 2.050 ;
        RECT  8.670 0.470 8.830 0.810 ;
        RECT  7.990 1.930 8.750 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  9.170 1.080 9.290 1.240 ;
        RECT  8.280 0.460 8.330 1.480 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  3.170 1.500 3.190 1.720 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
    END
END SEDFKCND1

MACRO SEDFKCND2
    CLASS CORE ;
    FOREIGN SEDFKCND2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.160 1.570 11.320 2.070 ;
        RECT  11.160 0.420 11.320 0.920 ;
        RECT  11.320 1.570 11.610 1.690 ;
        RECT  11.320 0.800 11.610 0.920 ;
        RECT  11.610 0.800 11.750 1.690 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 1.600 10.650 1.760 ;
        RECT  10.420 0.760 10.650 0.920 ;
        RECT  10.650 0.760 10.790 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.000 0.300 ;
        RECT  5.000 -0.300 5.220 0.340 ;
        RECT  5.220 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 5.230 2.820 ;
        RECT  5.230 2.180 5.450 2.820 ;
        RECT  5.450 2.220 5.830 2.820 ;
        RECT  5.830 2.180 6.050 2.820 ;
        RECT  6.050 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 9.350 2.820 ;
        RECT  9.350 2.180 9.570 2.820 ;
        RECT  9.570 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.330 0.460 8.440 1.740 ;
        RECT  8.440 1.360 8.490 1.740 ;
        RECT  8.490 1.360 9.745 1.480 ;
        RECT  9.745 1.090 9.905 1.480 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.310 1.740 ;
        RECT  3.310 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  10.170 1.080 10.530 1.240 ;
        RECT  10.050 0.710 10.170 1.760 ;
        RECT  9.560 0.710 10.050 0.870 ;
        RECT  9.730 1.600 10.050 1.760 ;
        RECT  9.440 0.710 9.560 1.240 ;
        RECT  11.040 1.080 11.290 1.240 ;
        RECT  10.920 0.470 11.040 2.050 ;
        RECT  9.250 0.470 10.920 0.590 ;
        RECT  8.970 1.930 10.920 2.050 ;
        RECT  9.090 0.470 9.250 0.690 ;
        RECT  8.830 0.570 9.090 0.690 ;
        RECT  8.750 1.630 8.970 2.050 ;
        RECT  8.670 0.570 8.830 0.810 ;
        RECT  7.990 1.930 8.750 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  9.170 1.080 9.440 1.240 ;
        RECT  8.280 0.460 8.330 1.480 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  3.170 1.500 3.190 1.740 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
    END
END SEDFKCND2

MACRO SEDFKCND4
    CLASS CORE ;
    FOREIGN SEDFKCND4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  12.110 1.650 12.430 2.030 ;
        RECT  12.110 0.490 12.430 0.870 ;
        RECT  12.430 0.490 12.850 2.030 ;
        RECT  12.850 1.650 13.020 2.030 ;
        RECT  12.850 0.490 13.020 0.870 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.710 1.600 11.150 1.760 ;
        RECT  10.710 0.760 11.150 0.920 ;
        RECT  11.150 0.760 11.570 1.760 ;
        RECT  11.570 1.600 11.660 1.760 ;
        RECT  11.570 0.760 11.660 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 13.440 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 8.930 2.820 ;
        RECT  8.930 2.180 9.150 2.820 ;
        RECT  9.150 2.220 13.440 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.310 1.740 ;
        RECT  3.310 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  8.440 1.150 10.150 1.300 ;
        RECT  8.400 1.670 8.540 1.810 ;
        RECT  8.400 0.460 8.440 1.300 ;
        RECT  10.460 1.080 10.840 1.240 ;
        RECT  10.340 0.710 10.460 1.810 ;
        RECT  9.850 0.710 10.340 0.870 ;
        RECT  10.020 1.650 10.340 1.810 ;
        RECT  9.730 0.710 9.850 1.030 ;
        RECT  11.940 1.080 12.215 1.240 ;
        RECT  11.820 0.470 11.940 2.050 ;
        RECT  9.540 0.470 11.820 0.590 ;
        RECT  9.550 1.930 11.820 2.050 ;
        RECT  9.330 1.930 9.550 2.090 ;
        RECT  9.380 0.470 9.540 0.690 ;
        RECT  8.830 0.570 9.380 0.690 ;
        RECT  8.870 1.930 9.330 2.050 ;
        RECT  8.710 1.620 8.870 2.050 ;
        RECT  8.670 0.570 8.830 0.810 ;
        RECT  7.990 1.930 8.710 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  9.320 0.890 9.730 1.030 ;
        RECT  8.280 0.460 8.400 1.810 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  3.170 1.500 3.190 1.740 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
        LAYER M1 ;
        RECT  12.110 1.650 12.215 2.030 ;
        RECT  12.110 0.490 12.215 0.870 ;
        RECT  10.710 1.600 10.935 1.760 ;
        RECT  10.710 0.760 10.935 0.920 ;
    END
END SEDFKCND4

MACRO SEDFKCNQD1
    CLASS CORE ;
    FOREIGN SEDFKCNQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.110 1.600 10.330 1.760 ;
        RECT  10.110 0.710 10.330 0.870 ;
        RECT  10.330 0.710 10.470 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.000 0.300 ;
        RECT  5.000 -0.300 5.220 0.340 ;
        RECT  5.220 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 10.510 0.300 ;
        RECT  10.510 -0.300 10.730 0.340 ;
        RECT  10.730 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 5.230 2.820 ;
        RECT  5.230 2.180 5.450 2.820 ;
        RECT  5.450 2.220 5.830 2.820 ;
        RECT  5.830 2.180 6.050 2.820 ;
        RECT  6.050 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 9.350 2.820 ;
        RECT  9.350 2.180 9.570 2.820 ;
        RECT  9.570 2.220 10.510 2.820 ;
        RECT  10.510 2.180 10.730 2.820 ;
        RECT  10.730 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.330 0.460 8.440 1.740 ;
        RECT  8.440 1.360 8.490 1.740 ;
        RECT  8.490 1.360 9.560 1.480 ;
        RECT  9.560 1.030 9.720 1.480 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.330 1.720 ;
        RECT  3.330 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  9.990 1.050 10.210 1.270 ;
        RECT  9.870 0.710 9.990 1.760 ;
        RECT  9.410 0.710 9.870 0.870 ;
        RECT  9.730 1.600 9.870 1.760 ;
        RECT  9.290 0.710 9.410 1.240 ;
        RECT  10.590 0.470 10.710 2.050 ;
        RECT  9.280 0.470 10.590 0.590 ;
        RECT  8.970 1.930 10.590 2.050 ;
        RECT  9.060 0.430 9.280 0.590 ;
        RECT  8.830 0.470 9.060 0.590 ;
        RECT  8.750 1.725 8.970 2.050 ;
        RECT  8.670 0.470 8.830 0.810 ;
        RECT  7.990 1.930 8.750 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  9.170 1.080 9.290 1.240 ;
        RECT  8.280 0.460 8.330 1.480 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  3.170 1.500 3.190 1.720 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
    END
END SEDFKCNQD1

MACRO SEDFKCNQD2
    CLASS CORE ;
    FOREIGN SEDFKCNQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.430 1.600 10.650 1.760 ;
        RECT  10.430 0.760 10.650 0.920 ;
        RECT  10.650 0.760 10.790 1.760 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.000 0.300 ;
        RECT  5.000 -0.300 5.220 0.340 ;
        RECT  5.220 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 10.850 0.300 ;
        RECT  10.850 -0.300 11.070 0.340 ;
        RECT  11.070 -0.300 11.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 5.230 2.820 ;
        RECT  5.230 2.180 5.450 2.820 ;
        RECT  5.450 2.220 5.830 2.820 ;
        RECT  5.830 2.180 6.050 2.820 ;
        RECT  6.050 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 9.350 2.820 ;
        RECT  9.350 2.180 9.570 2.820 ;
        RECT  9.570 2.220 10.850 2.820 ;
        RECT  10.850 2.180 11.070 2.820 ;
        RECT  11.070 2.220 11.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.330 0.460 8.440 1.740 ;
        RECT  8.440 1.360 8.490 1.740 ;
        RECT  8.490 1.360 9.745 1.480 ;
        RECT  9.745 1.090 9.905 1.480 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.310 1.740 ;
        RECT  3.310 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  10.170 1.080 10.530 1.240 ;
        RECT  10.050 0.710 10.170 1.760 ;
        RECT  9.560 0.710 10.050 0.870 ;
        RECT  9.730 1.600 10.050 1.760 ;
        RECT  9.440 0.710 9.560 1.240 ;
        RECT  10.920 0.470 11.040 2.050 ;
        RECT  9.250 0.470 10.920 0.590 ;
        RECT  8.970 1.930 10.920 2.050 ;
        RECT  9.090 0.470 9.250 0.690 ;
        RECT  8.830 0.570 9.090 0.690 ;
        RECT  8.750 1.720 8.970 2.050 ;
        RECT  8.670 0.570 8.830 0.810 ;
        RECT  7.990 1.930 8.750 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  9.170 1.080 9.440 1.240 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  8.280 0.460 8.330 1.480 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  3.170 1.500 3.190 1.740 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
    END
END SEDFKCNQD2

MACRO SEDFKCNQD4
    CLASS CORE ;
    FOREIGN SEDFKCNQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.840 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.285 4.070 1.515 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.005 4.710 1.570 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.420 1.600 10.830 1.760 ;
        RECT  10.420 0.760 10.830 0.920 ;
        RECT  10.830 0.760 11.250 1.760 ;
        RECT  11.250 1.600 11.370 1.760 ;
        RECT  11.250 0.760 11.370 0.920 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 0.725 0.250 1.250 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.050 1.005 1.510 1.235 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.670 1.235 ;
        END
    END CP
    PIN CN
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.470 1.235 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 3.550 0.300 ;
        RECT  3.550 -0.300 3.770 0.760 ;
        RECT  3.770 -0.300 5.660 0.300 ;
        RECT  5.660 -0.300 5.880 0.340 ;
        RECT  5.880 -0.300 7.450 0.300 ;
        RECT  7.450 -0.300 7.670 0.690 ;
        RECT  7.670 -0.300 11.840 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.450 2.820 ;
        RECT  0.450 1.690 0.670 2.820 ;
        RECT  0.670 2.220 1.750 2.820 ;
        RECT  1.750 2.180 1.970 2.820 ;
        RECT  1.970 2.220 2.390 2.820 ;
        RECT  2.390 2.180 2.610 2.820 ;
        RECT  2.610 2.220 3.670 2.820 ;
        RECT  3.670 2.030 3.890 2.820 ;
        RECT  3.890 2.220 7.530 2.820 ;
        RECT  7.530 2.030 7.750 2.820 ;
        RECT  7.750 2.220 9.350 2.820 ;
        RECT  9.350 2.180 9.570 2.820 ;
        RECT  9.570 2.220 11.840 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.440 1.150 9.860 1.300 ;
        RECT  7.480 0.810 7.900 0.930 ;
        RECT  7.900 1.510 8.020 1.670 ;
        RECT  7.900 0.560 8.020 0.930 ;
        RECT  8.020 0.560 8.060 1.670 ;
        RECT  8.060 0.810 8.140 1.670 ;
        RECT  7.000 0.610 7.160 1.750 ;
        RECT  7.160 1.270 7.730 1.390 ;
        RECT  7.730 1.050 7.890 1.390 ;
        RECT  6.060 0.710 6.350 0.870 ;
        RECT  6.350 0.710 6.470 1.570 ;
        RECT  6.470 1.100 6.880 1.260 ;
        RECT  6.590 1.400 6.810 1.810 ;
        RECT  4.390 0.470 6.420 0.590 ;
        RECT  6.420 0.430 6.660 0.590 ;
        RECT  5.240 0.710 5.820 0.870 ;
        RECT  5.820 0.710 5.940 1.570 ;
        RECT  5.940 1.080 6.200 1.240 ;
        RECT  4.830 1.410 4.940 1.570 ;
        RECT  4.580 0.710 4.940 0.870 ;
        RECT  4.940 0.710 5.060 1.570 ;
        RECT  3.190 0.780 3.310 1.740 ;
        RECT  3.310 0.780 3.350 1.030 ;
        RECT  3.350 0.910 4.210 1.030 ;
        RECT  4.210 0.910 4.370 1.560 ;
        RECT  2.840 0.470 2.880 0.910 ;
        RECT  2.880 0.470 3.000 1.810 ;
        RECT  3.000 0.470 3.290 0.630 ;
        RECT  1.590 1.360 1.710 1.840 ;
        RECT  1.710 1.360 1.740 1.480 ;
        RECT  1.410 0.710 1.740 0.850 ;
        RECT  1.740 0.710 1.860 1.480 ;
        RECT  1.860 1.360 2.130 1.480 ;
        RECT  2.130 1.360 2.290 1.810 ;
        RECT  2.290 1.360 2.600 1.480 ;
        RECT  2.600 1.095 2.760 1.480 ;
        RECT  0.920 0.470 2.150 0.590 ;
        RECT  2.150 0.470 2.310 0.710 ;
        RECT  0.260 1.380 0.460 1.500 ;
        RECT  0.070 0.440 0.460 0.600 ;
        RECT  0.460 0.440 0.580 1.500 ;
        RECT  0.580 1.330 0.800 1.500 ;
        RECT  0.800 1.360 1.470 1.500 ;
        RECT  8.400 1.670 8.540 1.810 ;
        RECT  8.400 0.460 8.440 1.300 ;
        RECT  10.170 1.080 10.550 1.240 ;
        RECT  10.050 0.710 10.170 1.810 ;
        RECT  9.560 0.710 10.050 0.870 ;
        RECT  9.730 1.650 10.050 1.810 ;
        RECT  9.440 0.710 9.560 1.030 ;
        RECT  11.530 0.470 11.650 2.050 ;
        RECT  9.250 0.470 11.530 0.590 ;
        RECT  8.870 1.930 11.530 2.050 ;
        RECT  9.090 0.470 9.250 0.690 ;
        RECT  8.830 0.570 9.090 0.690 ;
        RECT  8.710 1.660 8.870 2.050 ;
        RECT  8.670 0.570 8.830 0.810 ;
        RECT  7.990 1.930 8.710 2.050 ;
        RECT  7.870 1.790 7.990 2.050 ;
        RECT  7.410 1.790 7.870 1.910 ;
        RECT  7.290 1.790 7.410 2.050 ;
        RECT  4.130 1.930 7.290 2.050 ;
        RECT  4.010 1.790 4.130 2.050 ;
        RECT  3.550 1.790 4.010 1.910 ;
        RECT  3.430 1.790 3.550 2.050 ;
        RECT  2.010 1.930 3.430 2.050 ;
        RECT  9.170 0.890 9.440 1.030 ;
        RECT  8.280 0.460 8.400 1.810 ;
        RECT  7.320 0.810 7.480 1.080 ;
        RECT  6.780 0.610 7.000 0.770 ;
        RECT  6.210 1.410 6.350 1.570 ;
        RECT  4.320 1.690 6.590 1.810 ;
        RECT  4.230 0.470 4.390 0.790 ;
        RECT  5.460 1.410 5.820 1.570 ;
        RECT  3.170 1.500 3.190 1.740 ;
        RECT  1.850 1.600 2.010 2.050 ;
        RECT  2.820 1.590 2.880 1.810 ;
        RECT  1.060 1.680 1.590 1.840 ;
        RECT  0.760 0.470 0.920 0.710 ;
        RECT  0.100 1.380 0.260 1.900 ;
        LAYER M1 ;
        RECT  10.420 1.600 10.615 1.760 ;
        RECT  10.420 0.760 10.615 0.920 ;
    END
END SEDFKCNQD4

MACRO SEDFQD1
    CLASS CORE ;
    FOREIGN SEDFQD1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  9.660 1.580 9.690 1.800 ;
        RECT  9.660 0.720 9.690 0.940 ;
        RECT  9.690 0.720 9.830 1.800 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.350 ;
        RECT  6.110 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 10.030 0.300 ;
        RECT  10.030 -0.300 10.250 0.350 ;
        RECT  10.250 -0.300 10.880 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.730 2.820 ;
        RECT  5.730 2.170 5.950 2.820 ;
        RECT  5.950 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 8.990 2.820 ;
        RECT  8.990 2.170 9.210 2.820 ;
        RECT  9.210 2.220 10.030 2.820 ;
        RECT  10.030 2.170 10.250 2.820 ;
        RECT  10.250 2.220 10.880 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  7.380 1.810 7.955 1.930 ;
        RECT  7.955 1.810 8.075 2.050 ;
        RECT  8.075 1.930 10.530 2.050 ;
        RECT  10.410 1.520 10.530 1.680 ;
        RECT  10.410 0.730 10.530 0.890 ;
        RECT  10.530 0.730 10.650 2.050 ;
        RECT  8.830 0.800 9.390 0.960 ;
        RECT  9.300 0.420 9.390 0.590 ;
        RECT  9.390 0.420 9.510 1.800 ;
        RECT  9.510 0.420 9.540 0.590 ;
        RECT  9.540 0.470 10.150 0.590 ;
        RECT  10.150 0.470 10.270 1.280 ;
        RECT  10.270 1.060 10.410 1.280 ;
        RECT  8.580 0.420 8.700 1.270 ;
        RECT  8.270 1.670 8.960 1.810 ;
        RECT  8.700 1.140 8.960 1.270 ;
        RECT  8.960 1.140 9.080 1.810 ;
        RECT  9.080 1.140 9.270 1.360 ;
        RECT  8.410 1.390 8.720 1.550 ;
        RECT  7.540 1.440 8.020 1.600 ;
        RECT  7.990 0.530 8.020 0.770 ;
        RECT  8.020 0.530 8.140 1.600 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.560 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  9.270 1.640 9.390 1.800 ;
        RECT  8.320 0.420 8.580 0.560 ;
        RECT  8.260 0.790 8.410 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDFQD1

MACRO SEDFQD2
    CLASS CORE ;
    FOREIGN SEDFQD2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  10.010 0.750 10.150 1.770 ;
        RECT  10.150 1.610 10.350 1.770 ;
        RECT  10.150 0.750 10.350 0.910 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 5.890 0.300 ;
        RECT  5.890 -0.300 6.110 0.350 ;
        RECT  6.110 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 9.710 0.300 ;
        RECT  9.710 -0.300 9.930 0.340 ;
        RECT  9.930 -0.300 10.510 0.300 ;
        RECT  10.510 -0.300 10.730 0.350 ;
        RECT  10.730 -0.300 11.200 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 5.730 2.820 ;
        RECT  5.730 2.170 5.950 2.820 ;
        RECT  5.950 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 8.990 2.820 ;
        RECT  8.990 2.170 9.210 2.820 ;
        RECT  9.210 2.220 9.710 2.820 ;
        RECT  9.710 2.180 9.930 2.820 ;
        RECT  9.930 2.220 10.510 2.820 ;
        RECT  10.510 2.170 10.730 2.820 ;
        RECT  10.730 2.220 11.200 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  7.380 1.810 7.955 1.930 ;
        RECT  7.955 1.810 8.075 2.050 ;
        RECT  8.075 1.930 11.010 2.050 ;
        RECT  10.890 1.520 11.010 1.680 ;
        RECT  10.890 0.730 11.010 0.890 ;
        RECT  11.010 0.730 11.130 2.050 ;
        RECT  8.830 0.800 9.390 0.960 ;
        RECT  9.300 0.420 9.390 0.590 ;
        RECT  9.390 0.420 9.510 1.800 ;
        RECT  9.510 0.420 9.540 0.590 ;
        RECT  9.540 0.470 10.630 0.590 ;
        RECT  10.630 0.470 10.750 1.280 ;
        RECT  10.750 1.060 10.890 1.280 ;
        RECT  8.580 0.420 8.700 1.270 ;
        RECT  8.270 1.670 8.960 1.810 ;
        RECT  8.700 1.140 8.960 1.270 ;
        RECT  8.960 1.140 9.080 1.810 ;
        RECT  9.080 1.140 9.270 1.360 ;
        RECT  8.410 1.390 8.720 1.550 ;
        RECT  7.540 1.440 8.020 1.600 ;
        RECT  7.990 0.530 8.020 0.770 ;
        RECT  8.020 0.530 8.140 1.600 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.560 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  9.270 1.640 9.390 1.800 ;
        RECT  8.320 0.420 8.580 0.560 ;
        RECT  8.260 0.790 8.410 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
    END
END SEDFQD2

MACRO SEDFQD4
    CLASS CORE ;
    FOREIGN SEDFQD4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.610 1.005 3.850 1.235 ;
        RECT  3.850 1.005 4.010 1.450 ;
        RECT  4.010 1.005 4.070 1.235 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.530 0.890 4.690 1.130 ;
        RECT  4.690 0.890 4.890 1.010 ;
        RECT  4.890 0.445 5.030 1.010 ;
        END
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  11.110 1.520 11.470 1.680 ;
        RECT  11.110 0.750 11.470 0.910 ;
        RECT  11.470 0.750 11.890 1.680 ;
        RECT  11.890 1.520 12.060 1.680 ;
        RECT  11.890 0.750 12.060 0.910 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.070 0.730 1.290 ;
        RECT  0.730 1.070 0.870 1.810 ;
        RECT  0.870 1.690 0.900 1.810 ;
        RECT  0.900 1.690 1.020 1.840 ;
        RECT  1.020 1.720 1.340 1.840 ;
        RECT  1.340 1.720 1.460 1.910 ;
        RECT  1.460 1.790 1.910 1.910 ;
        RECT  1.910 1.790 2.040 2.050 ;
        RECT  2.040 1.930 2.470 2.050 ;
        RECT  2.470 1.930 2.710 2.100 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.370 1.285 1.700 1.515 ;
        RECT  1.700 1.080 1.830 1.515 ;
        RECT  1.830 1.080 1.890 1.300 ;
        END
    END D
    PIN CP
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 0.725 5.350 1.235 ;
        RECT  5.350 1.050 5.770 1.210 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 1.730 0.300 ;
        RECT  1.730 -0.300 1.950 0.460 ;
        RECT  1.950 -0.300 4.240 0.300 ;
        RECT  4.240 -0.300 4.460 0.510 ;
        RECT  4.460 -0.300 7.610 0.300 ;
        RECT  7.610 -0.300 7.770 0.770 ;
        RECT  7.770 -0.300 12.220 0.300 ;
        RECT  12.220 -0.300 12.440 0.340 ;
        RECT  12.440 -0.300 12.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 1.500 2.820 ;
        RECT  1.500 2.030 1.720 2.820 ;
        RECT  1.720 2.220 4.020 2.820 ;
        RECT  4.020 2.050 4.240 2.820 ;
        RECT  4.240 2.220 7.510 2.820 ;
        RECT  7.510 2.050 7.730 2.820 ;
        RECT  7.730 2.220 10.080 2.820 ;
        RECT  10.080 2.170 10.300 2.820 ;
        RECT  10.300 2.220 10.730 2.820 ;
        RECT  10.730 2.180 10.950 2.820 ;
        RECT  10.950 2.220 12.220 2.820 ;
        RECT  12.220 2.180 12.440 2.820 ;
        RECT  12.440 2.220 12.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  8.375 1.810 8.495 2.050 ;
        RECT  8.495 1.930 12.610 2.050 ;
        RECT  12.490 1.520 12.610 1.680 ;
        RECT  12.490 0.730 12.610 0.890 ;
        RECT  12.610 0.730 12.730 2.050 ;
        RECT  9.920 0.800 10.480 0.960 ;
        RECT  10.390 0.420 10.480 0.590 ;
        RECT  10.480 0.420 10.600 1.800 ;
        RECT  10.600 0.420 10.630 0.590 ;
        RECT  10.630 0.470 12.230 0.590 ;
        RECT  12.230 0.470 12.350 1.280 ;
        RECT  12.350 1.060 12.490 1.280 ;
        RECT  8.690 0.720 8.850 1.810 ;
        RECT  9.410 0.420 9.670 0.560 ;
        RECT  9.670 0.420 9.790 1.270 ;
        RECT  8.850 1.670 10.050 1.810 ;
        RECT  9.790 1.140 10.050 1.270 ;
        RECT  10.050 1.140 10.170 1.810 ;
        RECT  10.170 1.140 10.360 1.360 ;
        RECT  9.500 1.390 9.810 1.550 ;
        RECT  7.540 1.440 8.010 1.600 ;
        RECT  8.010 0.470 8.160 1.600 ;
        RECT  9.000 1.400 9.030 1.550 ;
        RECT  8.160 0.470 9.030 0.590 ;
        RECT  9.030 0.470 9.190 1.550 ;
        RECT  9.190 1.400 9.220 1.550 ;
        RECT  9.190 0.470 9.290 0.630 ;
        RECT  6.920 0.460 7.020 0.620 ;
        RECT  7.020 0.460 7.140 1.810 ;
        RECT  7.140 0.460 7.160 1.010 ;
        RECT  7.160 0.890 7.730 1.010 ;
        RECT  7.730 0.890 7.890 1.280 ;
        RECT  5.270 0.420 5.510 0.590 ;
        RECT  5.510 0.470 6.560 0.590 ;
        RECT  5.260 1.690 6.600 1.810 ;
        RECT  6.560 0.420 6.680 0.590 ;
        RECT  6.600 1.350 6.720 1.810 ;
        RECT  6.720 1.350 6.760 1.470 ;
        RECT  6.680 0.420 6.760 0.890 ;
        RECT  6.760 0.420 6.800 1.470 ;
        RECT  6.800 0.770 6.880 1.470 ;
        RECT  6.270 0.750 6.360 0.910 ;
        RECT  6.360 0.750 6.480 1.570 ;
        RECT  6.480 0.750 6.510 1.230 ;
        RECT  6.510 1.010 6.640 1.230 ;
        RECT  5.550 0.740 5.890 0.880 ;
        RECT  5.890 0.740 6.010 1.570 ;
        RECT  6.010 1.050 6.240 1.270 ;
        RECT  2.380 0.980 2.410 1.780 ;
        RECT  2.410 0.710 2.500 1.780 ;
        RECT  2.500 0.710 2.530 1.110 ;
        RECT  2.530 0.710 3.290 0.830 ;
        RECT  3.290 0.710 3.410 1.780 ;
        RECT  3.410 1.570 3.540 1.780 ;
        RECT  3.410 0.710 3.810 0.830 ;
        RECT  3.540 1.570 4.630 1.690 ;
        RECT  4.630 1.410 4.750 1.690 ;
        RECT  4.750 1.410 4.940 1.530 ;
        RECT  4.940 1.140 5.090 1.530 ;
        RECT  0.300 0.470 1.490 0.590 ;
        RECT  1.490 0.470 1.610 0.700 ;
        RECT  1.610 0.580 2.070 0.700 ;
        RECT  2.070 0.420 2.290 0.700 ;
        RECT  2.290 0.470 3.390 0.590 ;
        RECT  3.390 0.420 3.610 0.590 ;
        RECT  3.610 0.470 3.940 0.590 ;
        RECT  3.940 0.470 4.080 0.770 ;
        RECT  4.080 0.630 4.260 0.770 ;
        RECT  4.260 0.630 4.380 1.450 ;
        RECT  4.380 1.310 4.500 1.450 ;
        RECT  4.380 0.630 4.620 0.770 ;
        RECT  4.620 0.530 4.760 0.770 ;
        RECT  1.880 0.820 2.010 0.940 ;
        RECT  2.010 0.820 2.130 1.670 ;
        RECT  1.100 0.710 1.230 1.600 ;
        RECT  1.230 1.380 1.240 1.600 ;
        RECT  1.230 0.710 1.370 0.930 ;
        RECT  0.540 0.800 0.680 0.940 ;
        RECT  0.540 1.930 0.690 2.050 ;
        RECT  0.690 1.930 0.810 2.100 ;
        RECT  0.680 0.710 0.850 0.940 ;
        RECT  0.810 1.980 1.200 2.100 ;
        RECT  7.380 1.810 8.375 1.930 ;
        RECT  7.260 1.810 7.380 2.050 ;
        RECT  4.630 1.930 7.260 2.050 ;
        RECT  4.510 1.810 4.630 2.050 ;
        RECT  3.800 1.810 4.510 1.930 ;
        RECT  3.680 1.810 3.800 2.050 ;
        RECT  3.030 1.930 3.680 2.050 ;
        RECT  2.890 0.950 3.170 1.090 ;
        RECT  2.910 1.620 3.030 2.050 ;
        RECT  2.890 1.620 2.910 1.780 ;
        RECT  2.770 0.950 2.890 1.780 ;
        RECT  10.360 1.640 10.480 1.800 ;
        RECT  8.600 1.510 8.690 1.670 ;
        RECT  2.670 1.620 2.770 1.780 ;
        RECT  9.350 0.790 9.500 1.550 ;
        RECT  7.380 1.140 7.540 1.600 ;
        RECT  6.890 1.590 7.020 1.810 ;
        RECT  5.020 1.650 5.260 1.810 ;
        RECT  6.130 1.410 6.360 1.570 ;
        RECT  5.400 1.410 5.890 1.570 ;
        RECT  2.260 1.620 2.380 1.780 ;
        RECT  0.140 0.470 0.300 1.290 ;
        RECT  1.950 1.450 2.010 1.670 ;
        RECT  0.990 0.710 1.100 0.930 ;
        RECT  0.420 0.800 0.540 2.050 ;
        LAYER M1 ;
        RECT  11.110 0.750 11.255 0.910 ;
        RECT  11.110 1.520 11.255 1.680 ;
    END
END SEDFQD4

MACRO TIEH
    CLASS CORE ;
    FOREIGN TIEH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.960 0.390 2.100 ;
        RECT  0.390 1.005 0.550 2.100 ;
        RECT  0.550 1.960 0.580 2.100 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.360 0.420 0.580 0.870 ;
        RECT  0.240 0.750 0.360 0.870 ;
        RECT  0.080 0.750 0.240 1.290 ;
    END
END TIEH

MACRO TIEL
    CLASS CORE ;
    FOREIGN TIEL 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.640 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  0.390 0.420 0.550 1.235 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.640 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.640 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.550 1.960 0.580 2.100 ;
        RECT  0.390 1.390 0.550 2.100 ;
        RECT  0.240 1.390 0.390 1.510 ;
        RECT  0.080 1.030 0.240 1.510 ;
        RECT  0.360 1.960 0.390 2.100 ;
    END
END TIEL

MACRO XNR2D0
    CLASS CORE ;
    FOREIGN XNR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.490 2.790 1.900 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.510 0.300 ;
        RECT  0.510 -0.300 0.730 0.570 ;
        RECT  0.730 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.920 1.930 1.770 2.050 ;
        RECT  1.770 0.710 1.890 2.050 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.710 2.010 0.870 ;
        RECT  1.040 1.360 1.200 1.810 ;
        RECT  1.200 1.360 1.290 1.480 ;
        RECT  1.140 0.730 1.290 0.850 ;
        RECT  1.290 0.730 1.410 1.480 ;
        RECT  0.090 0.690 0.420 0.850 ;
        RECT  0.420 0.690 0.540 1.800 ;
        RECT  0.540 1.010 1.030 1.130 ;
        RECT  1.030 1.010 1.170 1.230 ;
        RECT  0.820 1.400 0.920 2.050 ;
        RECT  0.800 1.280 0.820 2.050 ;
        RECT  2.350 0.470 2.510 1.290 ;
        RECT  1.650 0.470 2.350 0.590 ;
        RECT  1.530 0.470 1.650 1.780 ;
        RECT  1.370 1.620 1.530 1.780 ;
        RECT  0.660 1.280 0.800 1.520 ;
        RECT  0.900 0.690 1.140 0.850 ;
        RECT  1.310 0.470 1.530 0.610 ;
        RECT  0.090 1.640 0.420 1.800 ;
    END
END XNR2D0

MACRO XNR2D1
    CLASS CORE ;
    FOREIGN XNR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.920 0.680 2.820 ;
        RECT  0.680 2.220 2.190 2.820 ;
        RECT  2.190 2.180 2.410 2.820 ;
        RECT  2.410 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.510 0.300 ;
        RECT  0.510 -0.300 0.730 0.570 ;
        RECT  0.730 -0.300 2.200 0.300 ;
        RECT  2.200 -0.300 2.420 0.340 ;
        RECT  2.420 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 1.260 0.820 2.050 ;
        RECT  0.820 1.380 0.920 2.050 ;
        RECT  0.920 1.930 1.770 2.050 ;
        RECT  1.770 0.710 1.890 2.050 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.710 2.010 0.870 ;
        RECT  1.040 1.360 1.200 1.810 ;
        RECT  1.200 1.360 1.290 1.480 ;
        RECT  1.140 0.730 1.290 0.850 ;
        RECT  1.290 0.730 1.410 1.480 ;
        RECT  0.090 0.690 0.420 0.850 ;
        RECT  0.420 0.690 0.540 1.800 ;
        RECT  0.540 1.010 1.030 1.130 ;
        RECT  1.030 1.010 1.170 1.230 ;
        RECT  2.350 0.470 2.510 1.290 ;
        RECT  1.650 0.470 2.350 0.590 ;
        RECT  1.530 0.470 1.650 1.780 ;
        RECT  1.310 0.470 1.530 0.610 ;
        RECT  1.370 1.620 1.530 1.780 ;
        RECT  0.660 1.260 0.800 1.500 ;
        RECT  0.900 0.690 1.140 0.850 ;
        RECT  0.090 1.640 0.420 1.800 ;
    END
END XNR2D1

MACRO XNR2D2
    CLASS CORE ;
    FOREIGN XNR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 1.960 2.865 2.100 ;
        RECT  2.865 1.390 2.970 2.100 ;
        RECT  2.865 0.420 2.970 0.900 ;
        RECT  2.970 0.420 3.025 2.100 ;
        RECT  3.025 1.960 3.055 2.100 ;
        RECT  3.025 0.780 3.110 1.515 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.285 1.050 2.310 1.270 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.530 2.820 ;
        RECT  0.530 2.180 0.750 2.820 ;
        RECT  0.750 2.220 2.445 2.820 ;
        RECT  2.445 2.180 2.665 2.820 ;
        RECT  2.665 2.220 3.520 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.530 0.300 ;
        RECT  0.530 -0.300 0.750 0.340 ;
        RECT  0.750 -0.300 3.520 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.275 0.470 1.395 0.850 ;
        RECT  1.315 1.360 1.475 1.810 ;
        RECT  1.395 0.680 1.495 0.850 ;
        RECT  1.475 1.360 1.565 1.480 ;
        RECT  1.495 0.730 1.565 0.850 ;
        RECT  1.565 0.730 1.685 1.480 ;
        RECT  0.905 0.710 1.025 0.870 ;
        RECT  1.025 0.710 1.145 1.800 ;
        RECT  1.145 1.010 1.445 1.230 ;
        RECT  0.305 0.470 1.275 0.590 ;
        RECT  2.165 0.710 2.365 0.870 ;
        RECT  2.165 1.640 2.285 1.800 ;
        RECT  2.045 0.710 2.165 2.050 ;
        RECT  0.565 1.930 2.045 2.050 ;
        RECT  2.745 1.050 2.805 1.270 ;
        RECT  2.625 0.470 2.745 1.270 ;
        RECT  1.925 0.470 2.625 0.590 ;
        RECT  1.805 0.470 1.925 1.780 ;
        RECT  1.665 0.470 1.805 0.610 ;
        RECT  1.645 1.620 1.805 1.780 ;
        RECT  0.425 1.020 0.565 2.050 ;
        RECT  0.145 0.470 0.305 1.975 ;
        RECT  0.905 1.640 1.025 1.800 ;
    END
END XNR2D2

MACRO XNR2D4
    CLASS CORE ;
    FOREIGN XNR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.420 1.650 4.750 2.030 ;
        RECT  4.420 0.490 4.750 0.870 ;
        RECT  4.750 0.490 5.170 2.030 ;
        RECT  5.170 1.650 5.330 2.030 ;
        RECT  5.170 0.490 5.330 0.870 ;
        END
    END ZN
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.600 1.005 3.760 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.150 0.710 3.160 0.850 ;
        RECT  2.310 0.950 2.690 1.080 ;
        RECT  2.690 0.950 2.810 1.330 ;
        RECT  2.810 1.180 2.910 1.330 ;
        RECT  1.420 0.470 1.560 0.630 ;
        RECT  1.560 0.470 1.680 1.810 ;
        RECT  1.680 0.470 2.220 0.590 ;
        RECT  1.680 1.690 2.440 1.810 ;
        RECT  2.220 0.430 2.460 0.590 ;
        RECT  3.030 0.710 3.150 2.050 ;
        RECT  2.920 0.710 3.030 0.850 ;
        RECT  2.990 1.570 3.030 2.050 ;
        RECT  0.970 1.930 2.990 2.050 ;
        RECT  0.940 1.080 1.440 1.240 ;
        RECT  0.940 1.930 0.970 2.100 ;
        RECT  0.780 0.420 0.940 2.100 ;
        RECT  0.750 1.930 0.780 2.100 ;
        RECT  0.280 1.930 0.750 2.050 ;
        RECT  0.250 1.930 0.280 2.100 ;
        RECT  0.090 0.420 0.250 2.100 ;
        RECT  3.420 0.710 3.960 0.870 ;
        RECT  3.420 1.640 3.920 1.800 ;
        RECT  3.300 0.710 3.420 1.800 ;
        RECT  4.280 1.080 4.530 1.240 ;
        RECT  4.160 0.470 4.280 2.040 ;
        RECT  3.540 0.470 4.160 0.590 ;
        RECT  3.560 1.920 4.160 2.040 ;
        RECT  3.320 1.920 3.560 2.080 ;
        RECT  3.320 0.430 3.540 0.590 ;
        RECT  2.750 0.470 3.320 0.590 ;
        RECT  2.580 1.450 2.820 1.610 ;
        RECT  2.590 0.470 2.750 0.830 ;
        RECT  1.950 0.710 2.590 0.830 ;
        RECT  2.040 1.450 2.580 1.570 ;
        RECT  1.950 1.430 2.040 1.570 ;
        RECT  1.820 0.710 1.950 1.570 ;
        RECT  3.270 1.150 3.300 1.370 ;
        RECT  0.060 1.960 0.090 2.100 ;
        RECT  2.070 0.950 2.310 1.100 ;
        RECT  1.420 1.670 1.560 1.810 ;
        LAYER M1 ;
        RECT  4.420 1.650 4.535 2.030 ;
        RECT  4.420 0.490 4.535 0.870 ;
    END
END XNR2D4

MACRO XNR3D0
    CLASS CORE ;
    FOREIGN XNR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.660 4.710 1.900 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.725 1.830 1.250 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.640 ;
        RECT  0.670 -0.300 1.920 0.300 ;
        RECT  1.920 -0.300 2.140 0.340 ;
        RECT  2.140 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.890 0.750 ;
        RECT  2.890 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.340 ;
        RECT  4.330 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.920 0.690 2.820 ;
        RECT  0.690 2.220 1.910 2.820 ;
        RECT  1.910 2.180 2.130 2.820 ;
        RECT  2.130 2.220 2.670 2.820 ;
        RECT  2.670 1.620 2.890 2.820 ;
        RECT  2.890 2.220 4.110 2.820 ;
        RECT  4.110 2.180 4.330 2.820 ;
        RECT  4.330 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.310 0.710 1.430 2.050 ;
        RECT  1.430 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.550 2.090 ;
        RECT  0.790 0.470 0.910 1.240 ;
        RECT  0.910 0.470 1.510 0.590 ;
        RECT  1.550 1.400 1.690 1.810 ;
        RECT  1.510 0.430 1.730 0.590 ;
        RECT  1.690 1.400 1.970 1.520 ;
        RECT  1.730 0.470 1.970 0.590 ;
        RECT  1.970 0.470 2.090 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.800 ;
        RECT  0.490 1.360 1.030 1.480 ;
        RECT  1.030 1.020 1.190 1.480 ;
        RECT  1.090 0.710 1.310 0.870 ;
        RECT  3.170 0.890 3.330 1.250 ;
        RECT  2.480 0.890 3.170 1.010 ;
        RECT  3.810 0.710 3.930 0.870 ;
        RECT  3.810 1.640 3.930 1.800 ;
        RECT  3.690 0.710 3.810 2.050 ;
        RECT  3.130 1.930 3.690 2.050 ;
        RECT  3.010 1.380 3.130 2.050 ;
        RECT  4.270 0.470 4.430 1.290 ;
        RECT  3.570 0.470 4.270 0.590 ;
        RECT  3.450 0.470 3.570 1.780 ;
        RECT  3.280 0.590 3.450 0.750 ;
        RECT  3.280 1.620 3.450 1.780 ;
        RECT  2.850 1.130 3.010 1.500 ;
        RECT  2.320 0.540 2.480 1.810 ;
        RECT  1.100 1.630 1.310 1.790 ;
        RECT  0.620 1.080 0.790 1.240 ;
        RECT  0.100 0.420 0.260 0.880 ;
    END
END XNR3D0

MACRO XNR3D1
    CLASS CORE ;
    FOREIGN XNR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.960 4.550 2.100 ;
        RECT  4.550 0.420 4.710 2.100 ;
        RECT  4.710 1.960 4.740 2.100 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.725 1.830 1.250 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.640 ;
        RECT  0.670 -0.300 1.920 0.300 ;
        RECT  1.920 -0.300 2.140 0.340 ;
        RECT  2.140 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.890 0.770 ;
        RECT  2.890 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.340 ;
        RECT  4.330 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.920 0.690 2.820 ;
        RECT  0.690 2.220 1.910 2.820 ;
        RECT  1.910 2.180 2.130 2.820 ;
        RECT  2.130 2.220 2.670 2.820 ;
        RECT  2.670 1.630 2.890 2.820 ;
        RECT  2.890 2.220 4.110 2.820 ;
        RECT  4.110 2.180 4.330 2.820 ;
        RECT  4.330 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.480 0.890 3.170 1.010 ;
        RECT  3.170 0.890 3.330 1.270 ;
        RECT  1.090 0.710 1.310 0.870 ;
        RECT  1.310 0.710 1.430 2.050 ;
        RECT  1.430 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.550 2.090 ;
        RECT  0.790 0.470 0.910 1.240 ;
        RECT  0.910 0.470 1.510 0.590 ;
        RECT  1.550 1.400 1.690 1.810 ;
        RECT  1.510 0.430 1.730 0.590 ;
        RECT  1.690 1.400 1.970 1.520 ;
        RECT  1.730 0.470 1.970 0.590 ;
        RECT  1.970 0.470 2.090 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.800 ;
        RECT  0.490 1.360 1.030 1.480 ;
        RECT  1.030 0.990 1.190 1.480 ;
        RECT  3.810 0.710 3.930 0.870 ;
        RECT  3.810 1.640 3.930 1.800 ;
        RECT  3.690 0.710 3.810 2.050 ;
        RECT  3.130 1.930 3.690 2.050 ;
        RECT  3.010 1.390 3.130 2.050 ;
        RECT  4.270 0.470 4.430 1.290 ;
        RECT  3.570 0.470 4.270 0.590 ;
        RECT  3.450 0.470 3.570 1.810 ;
        RECT  3.280 0.610 3.450 0.770 ;
        RECT  3.280 1.650 3.450 1.810 ;
        RECT  2.850 1.130 3.010 1.510 ;
        RECT  2.320 0.570 2.480 1.770 ;
        RECT  1.100 1.670 1.310 1.830 ;
        RECT  0.620 1.080 0.790 1.240 ;
        RECT  0.100 0.470 0.260 0.880 ;
    END
END XNR3D1

MACRO XNR3D2
    CLASS CORE ;
    FOREIGN XNR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.440 1.960 5.470 2.100 ;
        RECT  5.470 1.390 5.530 2.100 ;
        RECT  5.470 0.420 5.530 0.900 ;
        RECT  5.530 0.420 5.630 2.100 ;
        RECT  5.630 1.960 5.660 2.100 ;
        RECT  5.630 0.780 5.670 1.515 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.030 1.515 ;
        RECT  5.030 1.050 5.070 1.270 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.830 1.235 ;
        RECT  1.830 1.010 1.890 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.630 0.520 ;
        RECT  0.630 -0.300 2.710 0.300 ;
        RECT  2.710 -0.300 2.850 0.520 ;
        RECT  2.850 -0.300 6.080 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.710 2.820 ;
        RECT  2.710 1.980 2.850 2.820 ;
        RECT  2.850 2.220 6.080 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.970 0.470 3.090 0.760 ;
        RECT  3.090 0.470 3.370 0.590 ;
        RECT  3.370 0.420 3.590 0.590 ;
        RECT  1.440 1.690 1.745 1.810 ;
        RECT  1.745 1.690 1.865 2.050 ;
        RECT  1.865 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.570 2.090 ;
        RECT  0.970 0.470 1.640 0.590 ;
        RECT  1.620 1.400 1.860 1.570 ;
        RECT  1.640 0.430 1.860 0.590 ;
        RECT  1.860 1.400 2.030 1.520 ;
        RECT  1.860 0.470 2.030 0.590 ;
        RECT  2.030 0.470 2.150 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.910 ;
        RECT  0.490 1.790 0.915 1.910 ;
        RECT  0.915 1.790 1.035 2.050 ;
        RECT  1.035 1.930 1.380 2.050 ;
        RECT  1.380 1.930 1.620 2.090 ;
        RECT  2.480 0.640 2.970 0.760 ;
        RECT  3.950 0.720 4.090 1.810 ;
        RECT  3.350 1.690 3.950 1.810 ;
        RECT  4.770 0.710 4.920 0.870 ;
        RECT  4.770 1.715 4.910 1.875 ;
        RECT  4.650 0.710 4.770 2.050 ;
        RECT  3.090 1.930 4.650 2.050 ;
        RECT  2.970 1.050 3.090 2.050 ;
        RECT  5.350 1.050 5.390 1.290 ;
        RECT  5.230 0.470 5.350 1.290 ;
        RECT  4.470 0.470 5.230 0.590 ;
        RECT  4.310 0.470 4.470 1.670 ;
        RECT  3.830 0.470 4.310 0.590 ;
        RECT  3.710 0.470 3.830 1.570 ;
        RECT  3.520 0.760 3.710 0.920 ;
        RECT  3.520 1.430 3.710 1.570 ;
        RECT  2.930 1.050 2.970 1.290 ;
        RECT  3.210 0.710 3.350 1.810 ;
        RECT  2.320 0.640 2.480 1.710 ;
        RECT  1.280 0.720 1.440 1.810 ;
        RECT  0.750 0.420 0.970 0.590 ;
        RECT  0.100 0.640 0.260 0.880 ;
        RECT  0.900 0.710 1.060 1.670 ;
    END
END XNR3D2

MACRO XNR3D4
    CLASS CORE ;
    FOREIGN XNR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.650 6.990 2.030 ;
        RECT  6.670 0.490 6.990 0.870 ;
        RECT  6.990 0.490 7.410 2.030 ;
        RECT  7.410 1.650 7.580 2.030 ;
        RECT  7.410 0.490 7.580 0.870 ;
        END
    END ZN
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.620 0.520 ;
        RECT  0.620 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.050 1.690 2.170 2.050 ;
        RECT  2.170 1.930 3.410 2.050 ;
        RECT  3.410 1.930 3.630 2.090 ;
        RECT  3.630 1.930 4.730 2.050 ;
        RECT  4.730 1.930 4.950 2.090 ;
        RECT  2.850 1.450 3.030 1.570 ;
        RECT  2.850 0.550 3.100 0.710 ;
        RECT  3.100 0.470 3.220 0.710 ;
        RECT  3.030 1.450 3.250 1.670 ;
        RECT  3.220 0.470 4.020 0.590 ;
        RECT  3.250 1.450 4.050 1.570 ;
        RECT  0.960 0.470 1.620 0.590 ;
        RECT  1.620 0.430 1.840 0.590 ;
        RECT  1.600 1.430 2.310 1.570 ;
        RECT  1.840 0.470 2.310 0.590 ;
        RECT  2.310 1.430 2.410 1.810 ;
        RECT  2.310 0.470 2.410 0.890 ;
        RECT  2.410 0.470 2.530 1.810 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.250 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.910 ;
        RECT  0.490 1.790 0.895 1.910 ;
        RECT  0.895 1.790 1.015 2.050 ;
        RECT  1.015 1.930 1.410 2.050 ;
        RECT  1.410 1.930 1.650 2.090 ;
        RECT  1.420 1.690 2.050 1.810 ;
        RECT  4.670 1.190 4.970 1.310 ;
        RECT  4.670 1.450 4.790 1.570 ;
        RECT  4.550 1.190 4.670 1.570 ;
        RECT  3.280 1.210 4.550 1.330 ;
        RECT  5.410 0.710 6.220 0.870 ;
        RECT  5.980 1.410 6.200 1.810 ;
        RECT  5.410 1.410 5.980 1.570 ;
        RECT  5.280 0.710 5.410 1.570 ;
        RECT  4.430 0.950 5.280 1.070 ;
        RECT  4.310 0.950 4.430 1.090 ;
        RECT  6.530 1.080 6.775 1.240 ;
        RECT  6.410 0.470 6.530 2.050 ;
        RECT  5.130 0.470 6.410 0.590 ;
        RECT  5.190 1.930 6.410 2.050 ;
        RECT  5.070 1.650 5.190 2.050 ;
        RECT  4.910 0.430 5.130 0.590 ;
        RECT  4.910 1.650 5.070 1.810 ;
        RECT  4.340 0.470 4.910 0.590 ;
        RECT  3.390 1.690 4.910 1.810 ;
        RECT  4.220 0.470 4.340 0.830 ;
        RECT  3.390 0.710 4.220 0.830 ;
        RECT  3.890 0.970 4.310 1.090 ;
        RECT  4.470 0.710 4.970 0.830 ;
        RECT  3.140 0.880 3.280 1.330 ;
        RECT  1.260 0.720 1.420 1.810 ;
        RECT  2.730 0.550 2.850 1.570 ;
        RECT  0.740 0.420 0.960 0.590 ;
        RECT  0.090 0.640 0.250 0.880 ;
        RECT  0.880 0.710 1.040 1.670 ;
        LAYER M1 ;
        RECT  6.670 1.650 6.775 2.030 ;
        RECT  6.670 0.490 6.775 0.870 ;
    END
END XNR3D4

MACRO XNR4D0
    CLASS CORE ;
    FOREIGN XNR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 1.410 4.570 1.570 ;
        RECT  4.450 0.645 4.570 0.805 ;
        RECT  4.570 0.645 4.710 1.570 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.030 1.515 ;
        RECT  5.030 1.050 5.160 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 1.005 7.270 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 4.860 0.300 ;
        RECT  4.860 -0.300 5.080 0.340 ;
        RECT  5.080 -0.300 6.670 0.300 ;
        RECT  6.670 -0.300 6.890 0.530 ;
        RECT  6.890 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.820 2.820 ;
        RECT  2.820 1.960 3.040 2.820 ;
        RECT  3.040 2.220 4.870 2.820 ;
        RECT  4.870 2.180 5.090 2.820 ;
        RECT  5.090 2.220 6.670 2.820 ;
        RECT  6.670 2.030 6.890 2.820 ;
        RECT  6.890 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.720 1.610 3.880 1.770 ;
        RECT  3.000 1.070 3.120 1.230 ;
        RECT  6.070 0.710 6.190 0.850 ;
        RECT  5.230 1.410 5.280 1.570 ;
        RECT  5.950 1.160 6.070 1.860 ;
        RECT  6.070 1.740 6.870 1.860 ;
        RECT  6.870 0.650 6.990 1.860 ;
        RECT  6.990 1.700 7.290 1.860 ;
        RECT  6.990 0.650 7.290 0.810 ;
        RECT  5.280 0.470 5.450 1.570 ;
        RECT  5.450 0.470 6.430 0.590 ;
        RECT  6.430 0.470 6.550 1.240 ;
        RECT  6.550 1.080 6.670 1.240 ;
        RECT  6.190 0.710 6.310 1.620 ;
        RECT  6.310 1.480 6.430 1.620 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.150 0.590 ;
        RECT  4.150 0.470 4.310 1.810 ;
        RECT  4.310 1.690 5.630 1.810 ;
        RECT  5.630 0.720 5.750 1.810 ;
        RECT  5.750 1.590 5.820 1.810 ;
        RECT  5.750 0.720 5.870 0.860 ;
        RECT  3.880 1.610 3.900 2.050 ;
        RECT  3.720 0.710 3.900 0.850 ;
        RECT  3.900 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.300 2.050 ;
        RECT  4.300 1.930 4.540 2.090 ;
        RECT  2.620 1.690 3.205 1.810 ;
        RECT  3.205 1.690 3.325 2.050 ;
        RECT  3.325 1.890 3.720 2.050 ;
        RECT  3.360 0.710 3.460 0.850 ;
        RECT  3.460 0.710 3.580 1.570 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.480 2.050 ;
        RECT  2.480 1.930 2.700 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  2.460 0.590 2.620 1.810 ;
        RECT  3.330 1.430 3.460 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  5.910 1.160 5.950 1.400 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
    END
END XNR4D0

MACRO XNR4D1
    CLASS CORE ;
    FOREIGN XNR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 1.410 4.570 1.570 ;
        RECT  4.500 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.660 1.570 ;
        RECT  4.660 0.780 4.710 1.570 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.030 1.515 ;
        RECT  5.030 1.050 5.160 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 1.005 7.270 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 6.670 0.300 ;
        RECT  6.670 -0.300 6.890 0.530 ;
        RECT  6.890 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.820 2.820 ;
        RECT  2.820 1.960 3.040 2.820 ;
        RECT  3.040 2.220 6.670 2.820 ;
        RECT  6.670 2.030 6.890 2.820 ;
        RECT  6.890 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.190 0.710 6.310 1.620 ;
        RECT  6.310 1.480 6.430 1.620 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.150 0.590 ;
        RECT  4.150 0.470 4.310 1.810 ;
        RECT  6.550 1.080 6.670 1.240 ;
        RECT  4.310 1.690 5.630 1.810 ;
        RECT  5.630 0.720 5.750 1.810 ;
        RECT  5.750 1.590 5.820 1.810 ;
        RECT  5.750 0.720 5.870 0.860 ;
        RECT  3.880 1.610 3.900 2.050 ;
        RECT  3.720 0.710 3.900 0.850 ;
        RECT  3.900 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.300 2.050 ;
        RECT  4.300 1.930 4.540 2.090 ;
        RECT  2.620 1.690 3.205 1.810 ;
        RECT  3.205 1.690 3.325 2.050 ;
        RECT  3.325 1.890 3.720 2.050 ;
        RECT  3.360 0.710 3.460 0.850 ;
        RECT  6.430 0.470 6.550 1.240 ;
        RECT  3.460 0.710 3.580 1.570 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.480 2.050 ;
        RECT  2.480 1.930 2.700 2.090 ;
        RECT  5.450 0.470 6.430 0.590 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  5.280 0.470 5.450 1.570 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  6.990 0.650 7.290 0.810 ;
        RECT  6.990 1.700 7.290 1.860 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  6.870 0.650 6.990 1.860 ;
        RECT  6.070 1.740 6.870 1.860 ;
        RECT  5.950 1.160 6.070 1.860 ;
        RECT  5.910 1.160 5.950 1.400 ;
        RECT  5.230 1.410 5.280 1.570 ;
        RECT  6.070 0.710 6.190 0.850 ;
        RECT  3.000 1.070 3.120 1.230 ;
        RECT  3.720 1.610 3.880 1.770 ;
        RECT  2.460 0.590 2.620 1.810 ;
        RECT  3.330 1.430 3.460 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
    END
END XNR4D1

MACRO XNR4D2
    CLASS CORE ;
    FOREIGN XNR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.860 1.945 4.890 2.100 ;
        RECT  4.890 0.710 5.050 2.100 ;
        RECT  5.050 1.945 5.080 2.100 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.350 1.515 ;
        RECT  5.350 1.050 5.530 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 1.005 7.590 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.340 ;
        RECT  4.690 -0.300 7.020 0.300 ;
        RECT  7.020 -0.300 7.180 0.530 ;
        RECT  7.180 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.840 2.820 ;
        RECT  2.840 1.960 3.060 2.820 ;
        RECT  3.060 2.220 4.470 2.820 ;
        RECT  4.470 2.180 4.690 2.820 ;
        RECT  4.690 2.220 6.990 2.820 ;
        RECT  6.990 2.030 7.210 2.820 ;
        RECT  7.210 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.310 0.650 7.610 0.810 ;
        RECT  5.550 0.710 5.670 0.870 ;
        RECT  5.670 0.710 5.790 2.050 ;
        RECT  5.790 1.930 6.505 2.050 ;
        RECT  6.505 1.790 6.625 2.050 ;
        RECT  6.625 1.790 6.850 1.910 ;
        RECT  6.850 1.030 7.010 1.910 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.150 0.590 ;
        RECT  4.150 0.470 4.310 1.810 ;
        RECT  4.310 0.470 5.980 0.590 ;
        RECT  5.980 0.470 6.140 1.810 ;
        RECT  3.720 0.710 3.900 0.850 ;
        RECT  3.900 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.580 2.050 ;
        RECT  4.580 1.030 4.740 2.050 ;
        RECT  2.620 1.690 3.205 1.810 ;
        RECT  3.205 1.690 3.325 2.050 ;
        RECT  3.325 1.890 3.720 2.050 ;
        RECT  3.360 0.710 3.460 0.850 ;
        RECT  3.460 0.710 3.580 1.570 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.500 2.050 ;
        RECT  2.500 1.930 2.720 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  7.310 1.700 7.610 1.860 ;
        RECT  7.190 0.650 7.310 1.860 ;
        RECT  6.900 0.650 7.190 0.770 ;
        RECT  6.780 0.470 6.900 0.770 ;
        RECT  6.380 0.470 6.780 0.590 ;
        RECT  6.260 0.470 6.380 1.420 ;
        RECT  5.560 1.630 5.670 2.050 ;
        RECT  6.505 0.710 6.660 1.670 ;
        RECT  2.920 1.070 3.120 1.230 ;
        RECT  3.720 1.610 3.900 1.770 ;
        RECT  2.460 0.570 2.620 1.810 ;
        RECT  3.330 1.430 3.460 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
    END
END XNR4D2

MACRO XNR4D4
    CLASS CORE ;
    FOREIGN XNR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.320 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN ZN
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.800 1.650 5.070 2.030 ;
        RECT  4.780 0.760 5.070 0.920 ;
        RECT  5.070 0.760 5.490 2.030 ;
        RECT  5.490 1.650 5.720 2.030 ;
        RECT  5.490 0.760 5.740 0.920 ;
        END
    END ZN
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.850 1.005 5.990 1.515 ;
        RECT  5.990 1.050 6.170 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  8.070 1.005 8.230 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 7.660 0.300 ;
        RECT  7.660 -0.300 7.820 0.530 ;
        RECT  7.820 -0.300 8.320 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.840 2.820 ;
        RECT  2.840 1.960 3.060 2.820 ;
        RECT  3.060 2.220 7.630 2.820 ;
        RECT  7.630 2.030 7.850 2.820 ;
        RECT  7.850 2.220 8.320 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  6.310 0.710 6.430 2.050 ;
        RECT  6.430 1.930 7.145 2.050 ;
        RECT  7.145 1.790 7.265 2.050 ;
        RECT  7.265 1.790 7.490 1.910 ;
        RECT  7.490 1.030 7.650 1.910 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.150 0.590 ;
        RECT  4.150 0.470 4.310 1.810 ;
        RECT  4.310 0.470 6.620 0.590 ;
        RECT  6.620 0.470 6.780 1.810 ;
        RECT  3.720 0.710 3.900 0.850 ;
        RECT  3.900 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.520 2.050 ;
        RECT  4.520 1.030 4.680 2.050 ;
        RECT  2.620 1.690 3.205 1.810 ;
        RECT  3.205 1.690 3.325 2.050 ;
        RECT  3.325 1.890 3.720 2.050 ;
        RECT  3.360 0.710 3.460 0.850 ;
        RECT  3.460 0.710 3.580 1.570 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.500 2.050 ;
        RECT  2.500 1.930 2.720 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  6.190 0.710 6.310 0.870 ;
        RECT  7.950 0.650 8.250 0.810 ;
        RECT  7.950 1.700 8.250 1.860 ;
        RECT  7.830 0.650 7.950 1.860 ;
        RECT  7.540 0.650 7.830 0.770 ;
        RECT  7.420 0.470 7.540 0.770 ;
        RECT  7.020 0.470 7.420 0.590 ;
        RECT  6.900 0.470 7.020 1.420 ;
        RECT  6.200 1.630 6.310 2.050 ;
        RECT  7.145 0.710 7.300 1.670 ;
        RECT  2.920 1.070 3.120 1.230 ;
        RECT  3.720 1.610 3.900 1.770 ;
        RECT  2.460 0.570 2.620 1.810 ;
        RECT  3.330 1.430 3.460 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
        LAYER M1 ;
        RECT  5.705 1.650 5.720 2.030 ;
        RECT  5.705 0.760 5.740 0.920 ;
        RECT  4.800 1.650 4.855 2.030 ;
        RECT  4.780 0.760 4.855 0.920 ;
    END
END XNR4D4

MACRO XOR2D0
    CLASS CORE ;
    FOREIGN XOR2D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.630 0.610 2.790 1.840 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.030 2.190 1.510 ;
        RECT  2.190 1.390 2.330 1.510 ;
        RECT  2.330 1.390 2.470 2.075 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.990 1.040 1.235 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.590 2.820 ;
        RECT  0.590 1.560 0.810 2.820 ;
        RECT  0.810 2.220 2.230 2.820 ;
        RECT  2.230 2.200 2.450 2.820 ;
        RECT  2.450 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.420 0.300 ;
        RECT  0.420 -0.300 0.640 0.345 ;
        RECT  0.640 -0.300 2.230 0.300 ;
        RECT  2.230 -0.300 2.450 0.345 ;
        RECT  2.450 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.710 0.420 0.870 ;
        RECT  0.420 0.470 0.540 0.870 ;
        RECT  0.540 0.470 1.230 0.590 ;
        RECT  1.230 0.430 1.450 0.590 ;
        RECT  0.740 0.710 1.160 0.870 ;
        RECT  1.160 0.710 1.280 1.720 ;
        RECT  0.190 1.560 0.380 1.720 ;
        RECT  1.930 1.630 2.080 1.790 ;
        RECT  1.930 0.710 2.060 0.870 ;
        RECT  1.810 0.710 1.930 2.050 ;
        RECT  2.350 0.470 2.510 1.270 ;
        RECT  1.690 0.470 2.350 0.590 ;
        RECT  1.570 0.470 1.690 1.720 ;
        RECT  1.400 0.710 1.570 0.870 ;
        RECT  0.930 1.890 1.810 2.050 ;
        RECT  1.420 1.560 1.570 1.720 ;
        RECT  0.070 0.710 0.190 1.720 ;
        RECT  1.040 1.560 1.160 1.720 ;
    END
END XOR2D0

MACRO XOR2D1
    CLASS CORE ;
    FOREIGN XOR2D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.880 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.960 2.630 2.100 ;
        RECT  2.630 0.420 2.790 2.100 ;
        RECT  2.790 1.960 2.820 2.100 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.030 2.190 1.510 ;
        RECT  2.190 1.390 2.330 1.510 ;
        RECT  2.330 1.390 2.470 2.075 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.320 0.990 1.040 1.235 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.540 2.820 ;
        RECT  0.540 1.630 0.760 2.820 ;
        RECT  0.760 2.220 2.880 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.420 0.300 ;
        RECT  0.420 -0.300 0.640 0.345 ;
        RECT  0.640 -0.300 2.880 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.400 0.710 1.570 0.870 ;
        RECT  1.570 0.470 1.690 1.720 ;
        RECT  1.690 0.470 2.350 0.590 ;
        RECT  2.350 0.470 2.510 1.270 ;
        RECT  1.100 1.890 1.810 2.050 ;
        RECT  1.810 0.710 1.930 2.050 ;
        RECT  1.930 1.630 2.060 2.050 ;
        RECT  1.930 0.710 2.060 0.870 ;
        RECT  0.190 1.630 0.380 1.790 ;
        RECT  0.190 0.710 0.420 0.870 ;
        RECT  0.420 0.470 0.540 0.870 ;
        RECT  0.540 0.470 1.230 0.590 ;
        RECT  1.230 0.420 1.450 0.590 ;
        RECT  0.740 0.710 1.160 0.870 ;
        RECT  1.160 0.710 1.280 1.720 ;
        RECT  0.880 1.890 1.100 2.070 ;
        RECT  1.420 1.560 1.570 1.720 ;
        RECT  0.070 0.710 0.190 1.790 ;
        RECT  1.040 1.560 1.160 1.720 ;
    END
END XOR2D1

MACRO XOR2D2
    CLASS CORE ;
    FOREIGN XOR2D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.520 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  2.835 1.960 2.865 2.100 ;
        RECT  2.865 1.390 2.970 2.100 ;
        RECT  2.865 0.420 2.970 0.900 ;
        RECT  2.970 0.420 3.025 2.100 ;
        RECT  3.025 1.960 3.055 2.100 ;
        RECT  3.025 0.780 3.110 1.515 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.285 1.050 2.310 1.270 ;
        RECT  2.310 1.005 2.470 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.720 1.005 0.880 1.515 ;
        END
    END A1
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.530 2.820 ;
        RECT  0.530 2.180 0.750 2.820 ;
        RECT  0.750 2.220 2.445 2.820 ;
        RECT  2.445 2.180 2.665 2.820 ;
        RECT  2.665 2.220 3.520 2.820 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.530 0.300 ;
        RECT  0.530 -0.300 0.750 0.340 ;
        RECT  0.750 -0.300 3.520 0.300 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.275 0.470 1.395 0.850 ;
        RECT  1.315 1.360 1.475 1.810 ;
        RECT  1.395 0.640 1.495 0.850 ;
        RECT  1.475 1.360 1.565 1.480 ;
        RECT  1.495 0.730 1.565 0.850 ;
        RECT  1.565 0.730 1.685 1.480 ;
        RECT  0.905 0.710 1.025 0.870 ;
        RECT  1.025 0.710 1.145 1.800 ;
        RECT  1.145 1.060 1.405 1.220 ;
        RECT  0.305 0.470 1.275 0.590 ;
        RECT  2.165 0.710 2.365 0.870 ;
        RECT  2.165 1.640 2.285 1.800 ;
        RECT  2.045 0.710 2.165 2.050 ;
        RECT  0.565 1.930 2.045 2.050 ;
        RECT  2.745 1.050 2.805 1.270 ;
        RECT  2.625 0.470 2.745 1.270 ;
        RECT  1.925 0.470 2.625 0.590 ;
        RECT  1.805 0.470 1.925 1.780 ;
        RECT  1.665 0.470 1.805 0.610 ;
        RECT  1.645 1.620 1.805 1.780 ;
        RECT  0.425 1.020 0.565 2.050 ;
        RECT  0.145 0.470 0.305 1.960 ;
        RECT  0.905 1.640 1.025 1.800 ;
    END
END XOR2D2

MACRO XOR2D4
    CLASS CORE ;
    FOREIGN XOR2D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.430 1.650 4.750 2.030 ;
        RECT  4.430 0.490 4.750 0.870 ;
        RECT  4.750 0.490 5.170 2.030 ;
        RECT  5.170 1.650 5.340 2.030 ;
        RECT  5.170 0.490 5.340 0.870 ;
        END
    END Z
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.005 0.560 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.910 1.005 4.070 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.980 1.570 3.070 2.050 ;
        RECT  2.950 0.710 3.070 0.850 ;
        RECT  3.070 0.710 3.140 2.050 ;
        RECT  3.140 0.710 3.190 1.690 ;
        RECT  2.420 0.950 2.540 1.330 ;
        RECT  2.540 1.180 2.910 1.330 ;
        RECT  1.430 0.470 1.570 0.630 ;
        RECT  1.570 0.470 1.690 1.810 ;
        RECT  1.690 0.470 2.250 0.590 ;
        RECT  1.690 1.690 2.450 1.810 ;
        RECT  2.250 0.450 2.490 0.590 ;
        RECT  0.980 1.930 2.980 2.050 ;
        RECT  0.950 1.080 1.450 1.240 ;
        RECT  0.950 1.930 0.980 2.100 ;
        RECT  0.790 0.420 0.950 2.100 ;
        RECT  0.760 1.930 0.790 2.100 ;
        RECT  0.290 1.930 0.760 2.050 ;
        RECT  0.260 1.930 0.290 2.100 ;
        RECT  0.100 0.420 0.260 2.100 ;
        RECT  3.780 1.650 3.980 1.810 ;
        RECT  3.780 0.710 3.930 0.870 ;
        RECT  3.640 0.710 3.780 1.810 ;
        RECT  3.460 0.920 3.640 1.040 ;
        RECT  4.310 1.080 4.535 1.240 ;
        RECT  4.190 0.470 4.310 2.050 ;
        RECT  3.570 0.470 4.190 0.590 ;
        RECT  3.520 1.930 4.190 2.050 ;
        RECT  3.350 0.430 3.570 0.590 ;
        RECT  3.360 1.550 3.520 2.050 ;
        RECT  2.780 0.470 3.350 0.590 ;
        RECT  2.570 1.450 2.810 1.610 ;
        RECT  2.620 0.470 2.780 0.830 ;
        RECT  1.950 0.710 2.620 0.830 ;
        RECT  2.050 1.450 2.570 1.570 ;
        RECT  1.950 1.430 2.050 1.570 ;
        RECT  3.310 0.920 3.460 1.160 ;
        RECT  1.830 0.710 1.950 1.570 ;
        RECT  0.070 1.960 0.100 2.100 ;
        RECT  2.070 0.950 2.420 1.100 ;
        RECT  1.430 1.650 1.570 1.810 ;
        LAYER M1 ;
        RECT  4.430 1.650 4.535 2.030 ;
        RECT  4.430 0.490 4.535 0.870 ;
    END
END XOR2D4

MACRO XOR3D0
    CLASS CORE ;
    FOREIGN XOR3D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.550 0.660 4.710 1.900 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.725 1.830 1.250 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.640 ;
        RECT  0.670 -0.300 1.920 0.300 ;
        RECT  1.920 -0.300 2.140 0.340 ;
        RECT  2.140 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.890 0.750 ;
        RECT  2.890 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.340 ;
        RECT  4.330 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.920 0.690 2.820 ;
        RECT  0.690 2.220 1.910 2.820 ;
        RECT  1.910 2.180 2.130 2.820 ;
        RECT  2.130 2.220 2.670 2.820 ;
        RECT  2.670 1.620 2.890 2.820 ;
        RECT  2.890 2.220 4.110 2.820 ;
        RECT  4.110 2.180 4.330 2.820 ;
        RECT  4.330 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  1.310 0.710 1.430 2.050 ;
        RECT  1.430 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.550 2.090 ;
        RECT  0.790 0.470 0.910 1.240 ;
        RECT  0.910 0.470 1.510 0.590 ;
        RECT  1.550 1.400 1.690 1.810 ;
        RECT  1.510 0.430 1.730 0.590 ;
        RECT  1.690 1.400 1.970 1.520 ;
        RECT  1.730 0.470 1.970 0.590 ;
        RECT  1.970 0.470 2.090 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.800 ;
        RECT  0.490 1.360 1.030 1.480 ;
        RECT  1.030 1.160 1.190 1.480 ;
        RECT  1.090 0.710 1.310 0.870 ;
        RECT  3.170 0.890 3.330 1.250 ;
        RECT  2.480 0.890 3.170 1.010 ;
        RECT  3.810 0.710 3.930 0.870 ;
        RECT  3.810 1.640 3.930 1.800 ;
        RECT  3.690 0.710 3.810 2.050 ;
        RECT  3.130 1.930 3.690 2.050 ;
        RECT  3.010 1.380 3.130 2.050 ;
        RECT  4.270 0.470 4.430 1.290 ;
        RECT  3.570 0.470 4.270 0.590 ;
        RECT  3.450 0.470 3.570 1.780 ;
        RECT  3.280 1.620 3.450 1.780 ;
        RECT  3.280 0.590 3.450 0.750 ;
        RECT  2.850 1.130 3.010 1.500 ;
        RECT  2.320 0.540 2.480 1.810 ;
        RECT  1.100 1.630 1.310 1.790 ;
        RECT  0.620 1.080 0.790 1.240 ;
        RECT  0.100 0.420 0.260 0.880 ;
    END
END XOR3D0

MACRO XOR3D1
    CLASS CORE ;
    FOREIGN XOR3D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.960 4.550 2.100 ;
        RECT  4.550 0.420 4.710 2.100 ;
        RECT  4.710 1.960 4.740 2.100 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.005 4.090 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.670 0.725 1.830 1.250 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.450 0.300 ;
        RECT  0.450 -0.300 0.670 0.640 ;
        RECT  0.670 -0.300 1.920 0.300 ;
        RECT  1.920 -0.300 2.140 0.340 ;
        RECT  2.140 -0.300 2.670 0.300 ;
        RECT  2.670 -0.300 2.890 0.770 ;
        RECT  2.890 -0.300 4.110 0.300 ;
        RECT  4.110 -0.300 4.330 0.340 ;
        RECT  4.330 -0.300 4.800 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 1.920 0.690 2.820 ;
        RECT  0.690 2.220 1.910 2.820 ;
        RECT  1.910 2.180 2.130 2.820 ;
        RECT  2.130 2.220 2.670 2.820 ;
        RECT  2.670 1.630 2.890 2.820 ;
        RECT  2.890 2.220 4.110 2.820 ;
        RECT  4.110 2.180 4.330 2.820 ;
        RECT  4.330 2.220 4.800 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.810 0.710 3.930 0.870 ;
        RECT  2.480 0.890 3.170 1.010 ;
        RECT  3.170 0.890 3.330 1.270 ;
        RECT  1.090 0.710 1.310 0.870 ;
        RECT  1.310 0.710 1.430 2.050 ;
        RECT  1.430 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.550 2.090 ;
        RECT  0.790 0.470 0.910 1.240 ;
        RECT  0.910 0.470 1.510 0.590 ;
        RECT  1.550 1.400 1.690 1.810 ;
        RECT  1.510 0.430 1.730 0.590 ;
        RECT  1.690 1.400 1.970 1.520 ;
        RECT  1.730 0.470 1.970 0.590 ;
        RECT  1.970 0.470 2.090 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.800 ;
        RECT  0.490 1.360 1.030 1.480 ;
        RECT  1.030 1.170 1.190 1.480 ;
        RECT  3.810 1.640 3.930 1.800 ;
        RECT  3.690 0.710 3.810 2.050 ;
        RECT  3.130 1.930 3.690 2.050 ;
        RECT  3.010 1.390 3.130 2.050 ;
        RECT  4.270 0.470 4.430 1.290 ;
        RECT  3.570 0.470 4.270 0.590 ;
        RECT  3.450 0.470 3.570 1.810 ;
        RECT  3.280 0.610 3.450 0.770 ;
        RECT  2.850 1.130 3.010 1.510 ;
        RECT  3.280 1.650 3.450 1.810 ;
        RECT  2.320 0.570 2.480 1.770 ;
        RECT  1.100 1.700 1.310 1.860 ;
        RECT  0.620 1.080 0.790 1.240 ;
        RECT  0.100 0.470 0.260 0.880 ;
    END
END XOR3D1

MACRO XOR3D2
    CLASS CORE ;
    FOREIGN XOR3D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.760 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.710 1.410 4.890 1.550 ;
        RECT  4.760 0.420 4.890 0.900 ;
        RECT  4.890 0.420 4.920 1.550 ;
        RECT  4.920 0.780 5.030 1.550 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.170 1.050 4.250 1.270 ;
        RECT  4.250 1.005 4.390 1.790 ;
        RECT  4.390 1.670 5.260 1.790 ;
        RECT  5.260 1.030 5.420 1.790 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 0.725 1.830 1.235 ;
        RECT  1.830 1.010 1.900 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.490 0.300 ;
        RECT  0.490 -0.300 0.630 0.520 ;
        RECT  0.630 -0.300 2.040 0.300 ;
        RECT  2.040 -0.300 2.260 0.340 ;
        RECT  2.260 -0.300 2.710 0.300 ;
        RECT  2.710 -0.300 2.850 0.520 ;
        RECT  2.850 -0.300 4.330 0.300 ;
        RECT  4.330 -0.300 4.550 0.340 ;
        RECT  4.550 -0.300 5.760 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.710 2.820 ;
        RECT  2.710 1.980 2.850 2.820 ;
        RECT  2.850 2.220 4.330 2.820 ;
        RECT  4.330 2.180 4.550 2.820 ;
        RECT  4.550 2.220 5.760 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  5.500 0.440 5.570 0.940 ;
        RECT  5.570 0.440 5.660 2.050 ;
        RECT  5.660 0.820 5.690 2.050 ;
        RECT  3.730 0.470 4.520 0.590 ;
        RECT  4.520 0.470 4.640 1.270 ;
        RECT  4.640 1.050 4.770 1.270 ;
        RECT  2.480 0.640 2.970 0.760 ;
        RECT  2.970 0.470 3.090 0.760 ;
        RECT  3.090 0.470 3.250 0.590 ;
        RECT  3.250 0.420 3.470 0.590 ;
        RECT  1.280 0.720 1.440 1.830 ;
        RECT  1.440 1.680 1.470 1.830 ;
        RECT  1.470 1.710 1.745 1.830 ;
        RECT  1.745 1.710 1.865 2.050 ;
        RECT  1.865 1.930 2.330 2.050 ;
        RECT  2.330 1.930 2.570 2.090 ;
        RECT  0.970 0.470 1.640 0.590 ;
        RECT  1.620 1.400 1.860 1.570 ;
        RECT  1.640 0.430 1.860 0.590 ;
        RECT  1.860 1.400 2.080 1.520 ;
        RECT  1.860 0.470 2.080 0.590 ;
        RECT  2.080 0.470 2.200 1.520 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.260 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.910 ;
        RECT  0.490 1.790 0.915 1.910 ;
        RECT  0.915 1.790 1.035 2.100 ;
        RECT  1.035 1.980 1.290 2.100 ;
        RECT  4.030 1.910 5.570 2.050 ;
        RECT  4.030 0.710 4.180 0.870 ;
        RECT  3.910 0.710 4.030 2.050 ;
        RECT  3.090 1.930 3.910 2.050 ;
        RECT  2.970 1.050 3.090 2.050 ;
        RECT  2.930 1.050 2.970 1.290 ;
        RECT  3.590 0.470 3.730 1.680 ;
        RECT  2.320 0.640 2.480 1.770 ;
        RECT  3.210 0.720 3.350 1.680 ;
        RECT  1.250 1.680 1.280 1.830 ;
        RECT  0.750 0.420 0.970 0.590 ;
        RECT  0.100 0.640 0.260 0.880 ;
        RECT  0.900 0.710 1.060 1.670 ;
    END
END XOR3D2

MACRO XOR3D4
    CLASS CORE ;
    FOREIGN XOR3D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  6.670 1.650 6.990 2.030 ;
        RECT  6.670 0.490 6.990 0.870 ;
        RECT  6.990 0.490 7.410 2.030 ;
        RECT  7.410 1.650 7.580 2.030 ;
        RECT  7.410 0.490 7.580 0.870 ;
        END
    END Z
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.530 1.005 5.990 1.235 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.005 2.150 1.235 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.480 0.300 ;
        RECT  0.480 -0.300 0.620 0.520 ;
        RECT  0.620 -0.300 8.000 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.460 2.820 ;
        RECT  0.460 2.030 0.680 2.820 ;
        RECT  0.680 2.220 8.000 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.170 1.930 3.410 2.050 ;
        RECT  3.410 1.930 3.630 2.090 ;
        RECT  3.630 1.930 4.730 2.050 ;
        RECT  4.730 1.930 4.950 2.090 ;
        RECT  2.850 1.450 3.030 1.570 ;
        RECT  2.850 0.550 3.100 0.710 ;
        RECT  3.100 0.470 3.220 0.710 ;
        RECT  3.030 1.450 3.250 1.670 ;
        RECT  3.220 0.470 4.020 0.590 ;
        RECT  3.250 1.450 4.050 1.570 ;
        RECT  0.960 0.470 1.620 0.590 ;
        RECT  1.620 0.430 1.840 0.590 ;
        RECT  1.600 1.430 2.310 1.570 ;
        RECT  1.840 0.470 2.310 0.590 ;
        RECT  2.310 1.430 2.410 1.810 ;
        RECT  2.310 0.470 2.410 0.890 ;
        RECT  2.410 0.470 2.530 1.810 ;
        RECT  0.070 1.640 0.370 1.800 ;
        RECT  0.250 0.760 0.370 0.880 ;
        RECT  0.370 0.760 0.490 1.910 ;
        RECT  0.490 1.790 0.895 1.910 ;
        RECT  0.895 1.790 1.015 2.080 ;
        RECT  1.015 1.960 1.280 2.080 ;
        RECT  2.050 1.700 2.170 2.050 ;
        RECT  1.450 1.700 2.050 1.820 ;
        RECT  1.420 1.680 1.450 1.820 ;
        RECT  1.260 0.720 1.420 1.820 ;
        RECT  4.670 1.190 4.970 1.310 ;
        RECT  4.670 1.450 4.790 1.570 ;
        RECT  4.550 1.190 4.670 1.570 ;
        RECT  3.280 1.210 4.550 1.330 ;
        RECT  5.410 0.710 6.220 0.870 ;
        RECT  5.980 1.410 6.200 1.810 ;
        RECT  5.410 1.410 5.980 1.570 ;
        RECT  5.280 0.710 5.410 1.570 ;
        RECT  4.430 0.950 5.280 1.070 ;
        RECT  4.310 0.950 4.430 1.090 ;
        RECT  6.530 1.080 6.775 1.240 ;
        RECT  6.410 0.470 6.530 2.050 ;
        RECT  5.130 0.470 6.410 0.590 ;
        RECT  5.190 1.930 6.410 2.050 ;
        RECT  5.070 1.650 5.190 2.050 ;
        RECT  4.910 0.430 5.130 0.590 ;
        RECT  4.910 1.650 5.070 1.810 ;
        RECT  4.340 0.470 4.910 0.590 ;
        RECT  3.390 1.690 4.910 1.810 ;
        RECT  4.220 0.470 4.340 0.830 ;
        RECT  3.390 0.710 4.220 0.830 ;
        RECT  3.890 0.970 4.310 1.090 ;
        RECT  4.470 0.710 4.970 0.830 ;
        RECT  3.140 0.880 3.280 1.330 ;
        RECT  1.230 1.680 1.260 1.820 ;
        RECT  2.730 0.550 2.850 1.570 ;
        RECT  0.740 0.420 0.960 0.590 ;
        RECT  0.090 0.640 0.250 0.880 ;
        RECT  0.880 0.710 1.040 1.670 ;
        LAYER M1 ;
        RECT  6.670 1.650 6.775 2.030 ;
        RECT  6.670 0.490 6.775 0.870 ;
    END
END XOR3D4

MACRO XOR4D0
    CLASS CORE ;
    FOREIGN XOR4D0 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 1.410 4.570 1.570 ;
        RECT  4.450 0.645 4.570 0.805 ;
        RECT  4.570 0.645 4.710 1.570 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.030 1.515 ;
        RECT  5.030 1.050 5.160 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 1.005 7.270 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 4.860 0.300 ;
        RECT  4.860 -0.300 5.080 0.340 ;
        RECT  5.080 -0.300 6.670 0.300 ;
        RECT  6.670 -0.300 6.890 0.530 ;
        RECT  6.890 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.820 2.820 ;
        RECT  2.820 1.960 3.040 2.820 ;
        RECT  3.040 2.220 4.870 2.820 ;
        RECT  4.870 2.180 5.090 2.820 ;
        RECT  5.090 2.220 6.670 2.820 ;
        RECT  6.670 2.030 6.890 2.820 ;
        RECT  6.890 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.160 0.590 ;
        RECT  4.160 0.470 4.320 1.810 ;
        RECT  4.320 1.690 5.630 1.810 ;
        RECT  5.630 0.720 5.750 1.810 ;
        RECT  5.750 1.590 5.820 1.810 ;
        RECT  5.750 0.720 5.870 0.860 ;
        RECT  3.740 0.710 3.900 0.850 ;
        RECT  3.900 0.710 3.960 2.090 ;
        RECT  3.960 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.300 2.050 ;
        RECT  4.300 1.930 4.540 2.090 ;
        RECT  2.620 1.690 3.600 1.810 ;
        RECT  3.600 0.970 3.760 1.810 ;
        RECT  3.360 0.710 3.480 1.570 ;
        RECT  3.480 0.710 3.580 0.850 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.480 2.050 ;
        RECT  2.480 1.930 2.700 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  6.310 1.480 6.430 1.620 ;
        RECT  6.190 0.710 6.310 1.620 ;
        RECT  6.550 1.080 6.670 1.240 ;
        RECT  6.430 0.470 6.550 1.240 ;
        RECT  5.450 0.470 6.430 0.590 ;
        RECT  5.280 0.470 5.450 1.570 ;
        RECT  6.990 0.650 7.290 0.810 ;
        RECT  6.990 1.700 7.290 1.860 ;
        RECT  6.870 0.650 6.990 1.860 ;
        RECT  6.070 1.740 6.870 1.860 ;
        RECT  5.950 1.160 6.070 1.860 ;
        RECT  5.910 1.160 5.950 1.400 ;
        RECT  5.230 1.410 5.280 1.570 ;
        RECT  6.070 0.710 6.190 0.850 ;
        RECT  2.920 1.070 3.120 1.230 ;
        RECT  3.720 1.930 3.900 2.090 ;
        RECT  2.460 0.590 2.620 1.810 ;
        RECT  3.190 1.430 3.360 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
    END
END XOR4D0

MACRO XOR4D1
    CLASS CORE ;
    FOREIGN XOR4D1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.360 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.450 1.410 4.570 1.570 ;
        RECT  4.500 0.420 4.570 0.900 ;
        RECT  4.570 0.420 4.660 1.570 ;
        RECT  4.660 0.780 4.710 1.570 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  4.890 1.005 5.030 1.515 ;
        RECT  5.030 1.050 5.160 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.110 1.005 7.270 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 6.670 0.300 ;
        RECT  6.670 -0.300 6.890 0.530 ;
        RECT  6.890 -0.300 7.360 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.820 2.820 ;
        RECT  2.820 1.960 3.040 2.820 ;
        RECT  3.040 2.220 6.670 2.820 ;
        RECT  6.670 2.030 6.890 2.820 ;
        RECT  6.890 2.220 7.360 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  5.910 1.160 5.950 1.400 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  3.190 1.430 3.360 1.570 ;
        RECT  2.460 0.590 2.620 1.810 ;
        RECT  3.720 1.930 3.900 2.090 ;
        RECT  2.920 1.070 3.120 1.230 ;
        RECT  6.070 0.710 6.190 0.850 ;
        RECT  5.230 1.410 5.280 1.570 ;
        RECT  5.950 1.160 6.070 1.860 ;
        RECT  6.070 1.740 6.870 1.860 ;
        RECT  6.870 0.650 6.990 1.860 ;
        RECT  6.990 1.700 7.290 1.860 ;
        RECT  6.990 0.650 7.290 0.810 ;
        RECT  5.280 0.470 5.450 1.570 ;
        RECT  5.450 0.470 6.430 0.590 ;
        RECT  6.430 0.470 6.550 1.240 ;
        RECT  6.550 1.080 6.670 1.240 ;
        RECT  6.190 0.710 6.310 1.620 ;
        RECT  6.310 1.480 6.430 1.620 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.160 0.590 ;
        RECT  4.160 0.470 4.320 1.810 ;
        RECT  4.320 1.690 5.630 1.810 ;
        RECT  5.630 0.720 5.750 1.810 ;
        RECT  5.750 1.590 5.820 1.810 ;
        RECT  5.750 0.720 5.870 0.860 ;
        RECT  3.740 0.710 3.900 0.850 ;
        RECT  3.900 0.710 3.960 2.090 ;
        RECT  3.960 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.300 2.050 ;
        RECT  4.300 1.930 4.540 2.090 ;
        RECT  2.620 1.690 3.600 1.810 ;
        RECT  3.600 0.970 3.760 1.810 ;
        RECT  3.360 0.710 3.480 1.570 ;
        RECT  3.480 0.710 3.580 0.850 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.480 2.050 ;
        RECT  2.480 1.930 2.700 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  0.980 1.500 1.080 1.660 ;
    END
END XOR4D1

MACRO XOR4D2
    CLASS CORE ;
    FOREIGN XOR4D2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.680 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  4.860 1.945 4.890 2.100 ;
        RECT  4.890 0.710 5.050 2.100 ;
        RECT  5.050 1.945 5.080 2.100 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  5.210 1.005 5.350 1.515 ;
        RECT  5.350 1.050 5.530 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  7.430 1.005 7.590 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.180 0.300 ;
        RECT  2.180 -0.300 2.400 0.340 ;
        RECT  2.400 -0.300 2.840 0.300 ;
        RECT  2.840 -0.300 3.000 0.850 ;
        RECT  3.000 -0.300 4.470 0.300 ;
        RECT  4.470 -0.300 4.690 0.340 ;
        RECT  4.690 -0.300 7.020 0.300 ;
        RECT  7.020 -0.300 7.180 0.530 ;
        RECT  7.180 -0.300 7.680 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 2.170 2.820 ;
        RECT  2.170 2.180 2.390 2.820 ;
        RECT  2.390 2.220 2.820 2.820 ;
        RECT  2.820 1.960 3.040 2.820 ;
        RECT  3.040 2.220 4.470 2.820 ;
        RECT  4.470 2.180 4.690 2.820 ;
        RECT  4.690 2.220 6.990 2.820 ;
        RECT  6.990 2.030 7.210 2.820 ;
        RECT  7.210 2.220 7.680 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  7.310 1.700 7.610 1.860 ;
        RECT  7.310 0.650 7.610 0.810 ;
        RECT  5.550 0.710 5.670 0.870 ;
        RECT  5.670 0.710 5.790 2.050 ;
        RECT  5.790 1.930 6.505 2.050 ;
        RECT  6.505 1.790 6.625 2.050 ;
        RECT  6.625 1.790 6.850 1.910 ;
        RECT  6.850 1.030 7.010 1.910 ;
        RECT  3.120 0.470 3.240 1.230 ;
        RECT  3.240 0.470 4.160 0.590 ;
        RECT  4.160 0.470 4.320 1.810 ;
        RECT  4.320 0.470 5.980 0.590 ;
        RECT  5.980 0.470 6.140 1.810 ;
        RECT  3.720 0.710 3.900 0.850 ;
        RECT  3.900 0.710 3.960 2.090 ;
        RECT  3.960 0.710 4.020 2.050 ;
        RECT  4.020 1.930 4.580 2.050 ;
        RECT  4.580 1.030 4.740 2.050 ;
        RECT  2.620 1.690 3.600 1.810 ;
        RECT  3.600 1.005 3.760 1.810 ;
        RECT  3.360 0.710 3.480 1.570 ;
        RECT  3.480 0.710 3.600 0.850 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.480 2.050 ;
        RECT  2.480 1.930 2.700 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  7.190 0.650 7.310 1.860 ;
        RECT  6.900 0.650 7.190 0.770 ;
        RECT  6.780 0.470 6.900 0.770 ;
        RECT  6.380 0.470 6.780 0.590 ;
        RECT  5.560 1.630 5.670 2.050 ;
        RECT  6.505 0.710 6.660 1.670 ;
        RECT  2.920 1.070 3.120 1.230 ;
        RECT  3.720 1.930 3.900 2.090 ;
        RECT  2.460 0.570 2.620 1.810 ;
        RECT  3.240 1.430 3.360 1.570 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
        RECT  6.260 0.470 6.380 1.420 ;
    END
END XOR4D2

MACRO XOR4D4
    CLASS CORE ;
    FOREIGN XOR4D4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.280 BY 2.520 ;
    SYMMETRY x y ;
    SITE core ;
    PIN Z
        DIRECTION OUTPUT ;
        PORT
        LAYER M1 ;
        RECT  5.120 1.650 5.390 2.030 ;
        RECT  5.090 0.760 5.390 0.920 ;
        RECT  5.390 0.760 5.810 2.030 ;
        RECT  5.810 1.650 6.030 2.030 ;
        RECT  5.810 0.760 6.050 0.920 ;
        END
    END Z
    PIN A4
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  0.090 1.005 0.250 1.515 ;
        END
    END A4
    PIN A3
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  2.010 1.005 2.170 1.515 ;
        END
    END A3
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.005 6.950 1.515 ;
        RECT  6.950 1.050 7.120 1.270 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER M1 ;
        RECT  9.030 1.005 9.190 1.515 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.300 0.500 0.300 ;
        RECT  0.500 -0.300 0.640 0.570 ;
        RECT  0.640 -0.300 2.175 0.300 ;
        RECT  2.175 -0.300 2.395 0.340 ;
        RECT  2.395 -0.300 3.200 0.300 ;
        RECT  3.200 -0.300 3.420 0.340 ;
        RECT  3.420 -0.300 8.610 0.300 ;
        RECT  8.610 -0.300 8.770 0.530 ;
        RECT  8.770 -0.300 9.280 0.300 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 2.220 0.470 2.820 ;
        RECT  0.470 2.030 0.690 2.820 ;
        RECT  0.690 2.220 3.200 2.820 ;
        RECT  3.200 1.910 3.420 2.820 ;
        RECT  3.420 2.220 8.580 2.820 ;
        RECT  8.580 2.030 8.800 2.820 ;
        RECT  8.800 2.220 9.280 2.820 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  4.010 0.710 4.190 0.850 ;
        RECT  4.190 0.710 4.310 2.050 ;
        RECT  4.310 1.930 4.870 2.050 ;
        RECT  4.870 1.050 4.990 2.050 ;
        RECT  4.990 1.050 5.090 1.270 ;
        RECT  2.660 1.670 3.950 1.790 ;
        RECT  3.950 1.020 4.070 1.790 ;
        RECT  2.840 0.640 3.000 1.550 ;
        RECT  3.000 1.410 3.650 1.550 ;
        RECT  3.650 0.710 3.770 1.550 ;
        RECT  3.770 1.410 3.820 1.550 ;
        RECT  3.770 0.710 3.890 0.850 ;
        RECT  1.370 0.710 1.490 0.870 ;
        RECT  1.490 0.710 1.610 2.050 ;
        RECT  1.610 1.930 2.400 2.050 ;
        RECT  2.400 1.930 2.640 2.090 ;
        RECT  0.760 0.470 0.880 1.290 ;
        RECT  0.880 0.470 1.770 0.590 ;
        RECT  1.770 0.470 1.890 1.800 ;
        RECT  1.890 1.640 2.010 1.800 ;
        RECT  1.890 0.470 2.020 0.630 ;
        RECT  0.070 0.690 0.370 0.850 ;
        RECT  0.370 0.690 0.490 1.910 ;
        RECT  0.490 1.790 1.030 1.910 ;
        RECT  1.030 1.790 1.150 2.100 ;
        RECT  1.150 1.940 1.360 2.100 ;
        RECT  1.000 0.710 1.080 0.870 ;
        RECT  1.080 0.710 1.220 1.660 ;
        RECT  7.570 0.470 7.730 1.810 ;
        RECT  4.660 0.470 7.570 0.590 ;
        RECT  4.600 0.470 4.660 1.180 ;
        RECT  4.500 0.470 4.600 1.810 ;
        RECT  3.530 0.470 4.500 0.590 ;
        RECT  4.440 1.020 4.500 1.810 ;
        RECT  3.410 0.470 3.530 1.225 ;
        RECT  8.440 1.030 8.600 1.910 ;
        RECT  8.215 1.790 8.440 1.910 ;
        RECT  8.095 1.790 8.215 2.050 ;
        RECT  7.380 1.930 8.095 2.050 ;
        RECT  7.260 0.710 7.380 2.050 ;
        RECT  6.450 0.710 7.260 0.870 ;
        RECT  7.150 1.630 7.260 2.050 ;
        RECT  6.680 1.930 7.150 2.050 ;
        RECT  8.900 0.650 9.220 0.810 ;
        RECT  8.900 1.700 9.220 1.860 ;
        RECT  8.780 0.650 8.900 1.860 ;
        RECT  8.490 0.650 8.780 0.770 ;
        RECT  8.370 0.470 8.490 0.770 ;
        RECT  7.970 0.470 8.370 0.590 ;
        RECT  6.460 1.630 6.680 2.050 ;
        RECT  8.095 0.710 8.250 1.670 ;
        RECT  3.210 1.065 3.410 1.225 ;
        RECT  4.010 1.910 4.190 2.050 ;
        RECT  2.500 0.660 2.660 1.790 ;
        RECT  2.810 1.405 2.840 1.550 ;
        RECT  1.370 1.640 1.490 1.800 ;
        RECT  0.720 1.050 0.760 1.290 ;
        RECT  7.850 0.470 7.970 1.420 ;
        RECT  0.070 1.750 0.370 1.910 ;
        RECT  0.980 1.500 1.080 1.660 ;
        LAYER M1 ;
        RECT  6.025 1.650 6.030 2.030 ;
        RECT  6.025 0.760 6.050 0.920 ;
        RECT  5.120 1.650 5.175 2.030 ;
        RECT  5.090 0.760 5.175 0.920 ;
    END
END XOR4D4

END LIBRARY
